/*module XOR128(
  input  [127:0] io_data_in_1,
  input  [127:0] io_data_in_2,
  output [127:0] io_data_out
);
  assign io_data_out = io_data_in_1 ^ io_data_in_2; // @[XOR32.scala 18:31]
endmodule
module XOR8(
  input  [7:0] io_data_in_1,
  input  [7:0] io_data_in_2,
  output [7:0] io_data_out
);
  assign io_data_out = io_data_in_1 ^ io_data_in_2; // @[XOR32.scala 31:31]
endmodule
module G_func(
  input  [31:0] io_data_in,
  input  [7:0]  io_rc_in,
  output [31:0] io_data_out
);
  wire [7:0] io_data_out_a_io_data_in_1; // @[XOR32.scala 35:19]
  wire [7:0] io_data_out_a_io_data_in_2; // @[XOR32.scala 35:19]
  wire [7:0] io_data_out_a_io_data_out; // @[XOR32.scala 35:19]
  wire [7:0] _GEN_1 = 8'h1 == io_data_in[15:8] ? 8'h7c : 8'h63; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_2 = 8'h2 == io_data_in[15:8] ? 8'h77 : _GEN_1; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_3 = 8'h3 == io_data_in[15:8] ? 8'h7b : _GEN_2; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_4 = 8'h4 == io_data_in[15:8] ? 8'hf2 : _GEN_3; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_5 = 8'h5 == io_data_in[15:8] ? 8'h6b : _GEN_4; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_6 = 8'h6 == io_data_in[15:8] ? 8'h6f : _GEN_5; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_7 = 8'h7 == io_data_in[15:8] ? 8'hc5 : _GEN_6; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_8 = 8'h8 == io_data_in[15:8] ? 8'h30 : _GEN_7; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_9 = 8'h9 == io_data_in[15:8] ? 8'h1 : _GEN_8; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_10 = 8'ha == io_data_in[15:8] ? 8'h67 : _GEN_9; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_11 = 8'hb == io_data_in[15:8] ? 8'h2b : _GEN_10; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_12 = 8'hc == io_data_in[15:8] ? 8'hfe : _GEN_11; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_13 = 8'hd == io_data_in[15:8] ? 8'hd7 : _GEN_12; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_14 = 8'he == io_data_in[15:8] ? 8'hab : _GEN_13; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_15 = 8'hf == io_data_in[15:8] ? 8'h76 : _GEN_14; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_16 = 8'h10 == io_data_in[15:8] ? 8'hca : _GEN_15; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_17 = 8'h11 == io_data_in[15:8] ? 8'h82 : _GEN_16; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_18 = 8'h12 == io_data_in[15:8] ? 8'hc9 : _GEN_17; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_19 = 8'h13 == io_data_in[15:8] ? 8'h7d : _GEN_18; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_20 = 8'h14 == io_data_in[15:8] ? 8'hfa : _GEN_19; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_21 = 8'h15 == io_data_in[15:8] ? 8'h59 : _GEN_20; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_22 = 8'h16 == io_data_in[15:8] ? 8'h47 : _GEN_21; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_23 = 8'h17 == io_data_in[15:8] ? 8'hf0 : _GEN_22; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_24 = 8'h18 == io_data_in[15:8] ? 8'had : _GEN_23; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_25 = 8'h19 == io_data_in[15:8] ? 8'hd4 : _GEN_24; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_26 = 8'h1a == io_data_in[15:8] ? 8'ha2 : _GEN_25; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_27 = 8'h1b == io_data_in[15:8] ? 8'haf : _GEN_26; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_28 = 8'h1c == io_data_in[15:8] ? 8'h9c : _GEN_27; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_29 = 8'h1d == io_data_in[15:8] ? 8'ha4 : _GEN_28; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_30 = 8'h1e == io_data_in[15:8] ? 8'h72 : _GEN_29; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_31 = 8'h1f == io_data_in[15:8] ? 8'hc0 : _GEN_30; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_32 = 8'h20 == io_data_in[15:8] ? 8'hb7 : _GEN_31; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_33 = 8'h21 == io_data_in[15:8] ? 8'hfd : _GEN_32; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_34 = 8'h22 == io_data_in[15:8] ? 8'h93 : _GEN_33; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_35 = 8'h23 == io_data_in[15:8] ? 8'h26 : _GEN_34; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_36 = 8'h24 == io_data_in[15:8] ? 8'h36 : _GEN_35; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_37 = 8'h25 == io_data_in[15:8] ? 8'h3f : _GEN_36; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_38 = 8'h26 == io_data_in[15:8] ? 8'hf7 : _GEN_37; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_39 = 8'h27 == io_data_in[15:8] ? 8'hcc : _GEN_38; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_40 = 8'h28 == io_data_in[15:8] ? 8'h34 : _GEN_39; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_41 = 8'h29 == io_data_in[15:8] ? 8'ha5 : _GEN_40; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_42 = 8'h2a == io_data_in[15:8] ? 8'he5 : _GEN_41; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_43 = 8'h2b == io_data_in[15:8] ? 8'hf1 : _GEN_42; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_44 = 8'h2c == io_data_in[15:8] ? 8'h71 : _GEN_43; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_45 = 8'h2d == io_data_in[15:8] ? 8'hd8 : _GEN_44; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_46 = 8'h2e == io_data_in[15:8] ? 8'h31 : _GEN_45; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_47 = 8'h2f == io_data_in[15:8] ? 8'h15 : _GEN_46; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_48 = 8'h30 == io_data_in[15:8] ? 8'h4 : _GEN_47; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_49 = 8'h31 == io_data_in[15:8] ? 8'hc7 : _GEN_48; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_50 = 8'h32 == io_data_in[15:8] ? 8'h23 : _GEN_49; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_51 = 8'h33 == io_data_in[15:8] ? 8'hc3 : _GEN_50; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_52 = 8'h34 == io_data_in[15:8] ? 8'h18 : _GEN_51; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_53 = 8'h35 == io_data_in[15:8] ? 8'h96 : _GEN_52; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_54 = 8'h36 == io_data_in[15:8] ? 8'h5 : _GEN_53; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_55 = 8'h37 == io_data_in[15:8] ? 8'h9a : _GEN_54; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_56 = 8'h38 == io_data_in[15:8] ? 8'h7 : _GEN_55; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_57 = 8'h39 == io_data_in[15:8] ? 8'h12 : _GEN_56; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_58 = 8'h3a == io_data_in[15:8] ? 8'h80 : _GEN_57; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_59 = 8'h3b == io_data_in[15:8] ? 8'he2 : _GEN_58; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_60 = 8'h3c == io_data_in[15:8] ? 8'heb : _GEN_59; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_61 = 8'h3d == io_data_in[15:8] ? 8'h27 : _GEN_60; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_62 = 8'h3e == io_data_in[15:8] ? 8'hb2 : _GEN_61; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_63 = 8'h3f == io_data_in[15:8] ? 8'h75 : _GEN_62; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_64 = 8'h40 == io_data_in[15:8] ? 8'h9 : _GEN_63; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_65 = 8'h41 == io_data_in[15:8] ? 8'h83 : _GEN_64; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_66 = 8'h42 == io_data_in[15:8] ? 8'h2c : _GEN_65; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_67 = 8'h43 == io_data_in[15:8] ? 8'h1a : _GEN_66; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_68 = 8'h44 == io_data_in[15:8] ? 8'h1b : _GEN_67; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_69 = 8'h45 == io_data_in[15:8] ? 8'h6e : _GEN_68; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_70 = 8'h46 == io_data_in[15:8] ? 8'h5a : _GEN_69; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_71 = 8'h47 == io_data_in[15:8] ? 8'ha0 : _GEN_70; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_72 = 8'h48 == io_data_in[15:8] ? 8'h52 : _GEN_71; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_73 = 8'h49 == io_data_in[15:8] ? 8'h3b : _GEN_72; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_74 = 8'h4a == io_data_in[15:8] ? 8'hd6 : _GEN_73; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_75 = 8'h4b == io_data_in[15:8] ? 8'hb3 : _GEN_74; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_76 = 8'h4c == io_data_in[15:8] ? 8'h29 : _GEN_75; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_77 = 8'h4d == io_data_in[15:8] ? 8'he3 : _GEN_76; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_78 = 8'h4e == io_data_in[15:8] ? 8'h2f : _GEN_77; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_79 = 8'h4f == io_data_in[15:8] ? 8'h84 : _GEN_78; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_80 = 8'h50 == io_data_in[15:8] ? 8'h53 : _GEN_79; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_81 = 8'h51 == io_data_in[15:8] ? 8'hd1 : _GEN_80; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_82 = 8'h52 == io_data_in[15:8] ? 8'h0 : _GEN_81; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_83 = 8'h53 == io_data_in[15:8] ? 8'hed : _GEN_82; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_84 = 8'h54 == io_data_in[15:8] ? 8'h20 : _GEN_83; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_85 = 8'h55 == io_data_in[15:8] ? 8'hfc : _GEN_84; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_86 = 8'h56 == io_data_in[15:8] ? 8'hb1 : _GEN_85; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_87 = 8'h57 == io_data_in[15:8] ? 8'h5b : _GEN_86; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_88 = 8'h58 == io_data_in[15:8] ? 8'h6a : _GEN_87; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_89 = 8'h59 == io_data_in[15:8] ? 8'hcb : _GEN_88; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_90 = 8'h5a == io_data_in[15:8] ? 8'hbe : _GEN_89; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_91 = 8'h5b == io_data_in[15:8] ? 8'h39 : _GEN_90; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_92 = 8'h5c == io_data_in[15:8] ? 8'h4a : _GEN_91; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_93 = 8'h5d == io_data_in[15:8] ? 8'h4c : _GEN_92; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_94 = 8'h5e == io_data_in[15:8] ? 8'h58 : _GEN_93; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_95 = 8'h5f == io_data_in[15:8] ? 8'hcf : _GEN_94; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_96 = 8'h60 == io_data_in[15:8] ? 8'hd0 : _GEN_95; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_97 = 8'h61 == io_data_in[15:8] ? 8'hef : _GEN_96; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_98 = 8'h62 == io_data_in[15:8] ? 8'haa : _GEN_97; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_99 = 8'h63 == io_data_in[15:8] ? 8'hfb : _GEN_98; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_100 = 8'h64 == io_data_in[15:8] ? 8'h43 : _GEN_99; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_101 = 8'h65 == io_data_in[15:8] ? 8'h4d : _GEN_100; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_102 = 8'h66 == io_data_in[15:8] ? 8'h33 : _GEN_101; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_103 = 8'h67 == io_data_in[15:8] ? 8'h85 : _GEN_102; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_104 = 8'h68 == io_data_in[15:8] ? 8'h45 : _GEN_103; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_105 = 8'h69 == io_data_in[15:8] ? 8'hf9 : _GEN_104; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_106 = 8'h6a == io_data_in[15:8] ? 8'h2 : _GEN_105; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_107 = 8'h6b == io_data_in[15:8] ? 8'h7f : _GEN_106; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_108 = 8'h6c == io_data_in[15:8] ? 8'h50 : _GEN_107; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_109 = 8'h6d == io_data_in[15:8] ? 8'h3c : _GEN_108; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_110 = 8'h6e == io_data_in[15:8] ? 8'h9f : _GEN_109; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_111 = 8'h6f == io_data_in[15:8] ? 8'ha8 : _GEN_110; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_112 = 8'h70 == io_data_in[15:8] ? 8'h51 : _GEN_111; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_113 = 8'h71 == io_data_in[15:8] ? 8'ha3 : _GEN_112; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_114 = 8'h72 == io_data_in[15:8] ? 8'h40 : _GEN_113; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_115 = 8'h73 == io_data_in[15:8] ? 8'h8f : _GEN_114; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_116 = 8'h74 == io_data_in[15:8] ? 8'h92 : _GEN_115; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_117 = 8'h75 == io_data_in[15:8] ? 8'h9d : _GEN_116; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_118 = 8'h76 == io_data_in[15:8] ? 8'h38 : _GEN_117; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_119 = 8'h77 == io_data_in[15:8] ? 8'hf5 : _GEN_118; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_120 = 8'h78 == io_data_in[15:8] ? 8'hbc : _GEN_119; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_121 = 8'h79 == io_data_in[15:8] ? 8'hb6 : _GEN_120; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_122 = 8'h7a == io_data_in[15:8] ? 8'hda : _GEN_121; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_123 = 8'h7b == io_data_in[15:8] ? 8'h21 : _GEN_122; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_124 = 8'h7c == io_data_in[15:8] ? 8'h10 : _GEN_123; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_125 = 8'h7d == io_data_in[15:8] ? 8'hff : _GEN_124; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_126 = 8'h7e == io_data_in[15:8] ? 8'hf3 : _GEN_125; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_127 = 8'h7f == io_data_in[15:8] ? 8'hd2 : _GEN_126; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_128 = 8'h80 == io_data_in[15:8] ? 8'hcd : _GEN_127; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_129 = 8'h81 == io_data_in[15:8] ? 8'hc : _GEN_128; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_130 = 8'h82 == io_data_in[15:8] ? 8'h13 : _GEN_129; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_131 = 8'h83 == io_data_in[15:8] ? 8'hec : _GEN_130; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_132 = 8'h84 == io_data_in[15:8] ? 8'h5f : _GEN_131; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_133 = 8'h85 == io_data_in[15:8] ? 8'h97 : _GEN_132; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_134 = 8'h86 == io_data_in[15:8] ? 8'h44 : _GEN_133; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_135 = 8'h87 == io_data_in[15:8] ? 8'h17 : _GEN_134; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_136 = 8'h88 == io_data_in[15:8] ? 8'hc4 : _GEN_135; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_137 = 8'h89 == io_data_in[15:8] ? 8'ha7 : _GEN_136; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_138 = 8'h8a == io_data_in[15:8] ? 8'h7e : _GEN_137; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_139 = 8'h8b == io_data_in[15:8] ? 8'h3d : _GEN_138; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_140 = 8'h8c == io_data_in[15:8] ? 8'h64 : _GEN_139; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_141 = 8'h8d == io_data_in[15:8] ? 8'h5d : _GEN_140; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_142 = 8'h8e == io_data_in[15:8] ? 8'h19 : _GEN_141; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_143 = 8'h8f == io_data_in[15:8] ? 8'h73 : _GEN_142; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_144 = 8'h90 == io_data_in[15:8] ? 8'h60 : _GEN_143; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_145 = 8'h91 == io_data_in[15:8] ? 8'h81 : _GEN_144; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_146 = 8'h92 == io_data_in[15:8] ? 8'h4f : _GEN_145; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_147 = 8'h93 == io_data_in[15:8] ? 8'hdc : _GEN_146; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_148 = 8'h94 == io_data_in[15:8] ? 8'h22 : _GEN_147; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_149 = 8'h95 == io_data_in[15:8] ? 8'h2a : _GEN_148; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_150 = 8'h96 == io_data_in[15:8] ? 8'h90 : _GEN_149; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_151 = 8'h97 == io_data_in[15:8] ? 8'h88 : _GEN_150; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_152 = 8'h98 == io_data_in[15:8] ? 8'h46 : _GEN_151; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_153 = 8'h99 == io_data_in[15:8] ? 8'hee : _GEN_152; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_154 = 8'h9a == io_data_in[15:8] ? 8'hb8 : _GEN_153; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_155 = 8'h9b == io_data_in[15:8] ? 8'h14 : _GEN_154; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_156 = 8'h9c == io_data_in[15:8] ? 8'hde : _GEN_155; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_157 = 8'h9d == io_data_in[15:8] ? 8'h5e : _GEN_156; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_158 = 8'h9e == io_data_in[15:8] ? 8'hb : _GEN_157; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_159 = 8'h9f == io_data_in[15:8] ? 8'hdb : _GEN_158; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_160 = 8'ha0 == io_data_in[15:8] ? 8'he0 : _GEN_159; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_161 = 8'ha1 == io_data_in[15:8] ? 8'h32 : _GEN_160; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_162 = 8'ha2 == io_data_in[15:8] ? 8'h3a : _GEN_161; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_163 = 8'ha3 == io_data_in[15:8] ? 8'ha : _GEN_162; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_164 = 8'ha4 == io_data_in[15:8] ? 8'h49 : _GEN_163; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_165 = 8'ha5 == io_data_in[15:8] ? 8'h6 : _GEN_164; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_166 = 8'ha6 == io_data_in[15:8] ? 8'h24 : _GEN_165; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_167 = 8'ha7 == io_data_in[15:8] ? 8'h5c : _GEN_166; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_168 = 8'ha8 == io_data_in[15:8] ? 8'hc2 : _GEN_167; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_169 = 8'ha9 == io_data_in[15:8] ? 8'hd3 : _GEN_168; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_170 = 8'haa == io_data_in[15:8] ? 8'hac : _GEN_169; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_171 = 8'hab == io_data_in[15:8] ? 8'h62 : _GEN_170; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_172 = 8'hac == io_data_in[15:8] ? 8'h91 : _GEN_171; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_173 = 8'had == io_data_in[15:8] ? 8'h95 : _GEN_172; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_174 = 8'hae == io_data_in[15:8] ? 8'he4 : _GEN_173; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_175 = 8'haf == io_data_in[15:8] ? 8'h79 : _GEN_174; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_176 = 8'hb0 == io_data_in[15:8] ? 8'he7 : _GEN_175; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_177 = 8'hb1 == io_data_in[15:8] ? 8'hc8 : _GEN_176; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_178 = 8'hb2 == io_data_in[15:8] ? 8'h37 : _GEN_177; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_179 = 8'hb3 == io_data_in[15:8] ? 8'h6d : _GEN_178; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_180 = 8'hb4 == io_data_in[15:8] ? 8'h8d : _GEN_179; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_181 = 8'hb5 == io_data_in[15:8] ? 8'hd5 : _GEN_180; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_182 = 8'hb6 == io_data_in[15:8] ? 8'h4e : _GEN_181; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_183 = 8'hb7 == io_data_in[15:8] ? 8'ha9 : _GEN_182; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_184 = 8'hb8 == io_data_in[15:8] ? 8'h6c : _GEN_183; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_185 = 8'hb9 == io_data_in[15:8] ? 8'h56 : _GEN_184; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_186 = 8'hba == io_data_in[15:8] ? 8'hf4 : _GEN_185; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_187 = 8'hbb == io_data_in[15:8] ? 8'hea : _GEN_186; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_188 = 8'hbc == io_data_in[15:8] ? 8'h65 : _GEN_187; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_189 = 8'hbd == io_data_in[15:8] ? 8'h7a : _GEN_188; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_190 = 8'hbe == io_data_in[15:8] ? 8'hae : _GEN_189; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_191 = 8'hbf == io_data_in[15:8] ? 8'h8 : _GEN_190; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_192 = 8'hc0 == io_data_in[15:8] ? 8'hba : _GEN_191; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_193 = 8'hc1 == io_data_in[15:8] ? 8'h78 : _GEN_192; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_194 = 8'hc2 == io_data_in[15:8] ? 8'h25 : _GEN_193; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_195 = 8'hc3 == io_data_in[15:8] ? 8'h2e : _GEN_194; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_196 = 8'hc4 == io_data_in[15:8] ? 8'h1c : _GEN_195; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_197 = 8'hc5 == io_data_in[15:8] ? 8'ha6 : _GEN_196; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_198 = 8'hc6 == io_data_in[15:8] ? 8'hb4 : _GEN_197; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_199 = 8'hc7 == io_data_in[15:8] ? 8'hc6 : _GEN_198; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_200 = 8'hc8 == io_data_in[15:8] ? 8'he8 : _GEN_199; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_201 = 8'hc9 == io_data_in[15:8] ? 8'hdd : _GEN_200; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_202 = 8'hca == io_data_in[15:8] ? 8'h74 : _GEN_201; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_203 = 8'hcb == io_data_in[15:8] ? 8'h1f : _GEN_202; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_204 = 8'hcc == io_data_in[15:8] ? 8'h4b : _GEN_203; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_205 = 8'hcd == io_data_in[15:8] ? 8'hbd : _GEN_204; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_206 = 8'hce == io_data_in[15:8] ? 8'h8b : _GEN_205; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_207 = 8'hcf == io_data_in[15:8] ? 8'h8a : _GEN_206; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_208 = 8'hd0 == io_data_in[15:8] ? 8'h70 : _GEN_207; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_209 = 8'hd1 == io_data_in[15:8] ? 8'h3e : _GEN_208; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_210 = 8'hd2 == io_data_in[15:8] ? 8'hb5 : _GEN_209; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_211 = 8'hd3 == io_data_in[15:8] ? 8'h66 : _GEN_210; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_212 = 8'hd4 == io_data_in[15:8] ? 8'h48 : _GEN_211; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_213 = 8'hd5 == io_data_in[15:8] ? 8'h3 : _GEN_212; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_214 = 8'hd6 == io_data_in[15:8] ? 8'hf6 : _GEN_213; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_215 = 8'hd7 == io_data_in[15:8] ? 8'he : _GEN_214; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_216 = 8'hd8 == io_data_in[15:8] ? 8'h61 : _GEN_215; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_217 = 8'hd9 == io_data_in[15:8] ? 8'h35 : _GEN_216; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_218 = 8'hda == io_data_in[15:8] ? 8'h57 : _GEN_217; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_219 = 8'hdb == io_data_in[15:8] ? 8'hb9 : _GEN_218; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_220 = 8'hdc == io_data_in[15:8] ? 8'h86 : _GEN_219; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_221 = 8'hdd == io_data_in[15:8] ? 8'hc1 : _GEN_220; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_222 = 8'hde == io_data_in[15:8] ? 8'h1d : _GEN_221; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_223 = 8'hdf == io_data_in[15:8] ? 8'h9e : _GEN_222; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_224 = 8'he0 == io_data_in[15:8] ? 8'he1 : _GEN_223; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_225 = 8'he1 == io_data_in[15:8] ? 8'hf8 : _GEN_224; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_226 = 8'he2 == io_data_in[15:8] ? 8'h98 : _GEN_225; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_227 = 8'he3 == io_data_in[15:8] ? 8'h11 : _GEN_226; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_228 = 8'he4 == io_data_in[15:8] ? 8'h69 : _GEN_227; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_229 = 8'he5 == io_data_in[15:8] ? 8'hd9 : _GEN_228; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_230 = 8'he6 == io_data_in[15:8] ? 8'h8e : _GEN_229; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_231 = 8'he7 == io_data_in[15:8] ? 8'h94 : _GEN_230; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_232 = 8'he8 == io_data_in[15:8] ? 8'h9b : _GEN_231; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_233 = 8'he9 == io_data_in[15:8] ? 8'h1e : _GEN_232; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_234 = 8'hea == io_data_in[15:8] ? 8'h87 : _GEN_233; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_235 = 8'heb == io_data_in[15:8] ? 8'he9 : _GEN_234; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_236 = 8'hec == io_data_in[15:8] ? 8'hce : _GEN_235; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_237 = 8'hed == io_data_in[15:8] ? 8'h55 : _GEN_236; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_238 = 8'hee == io_data_in[15:8] ? 8'h28 : _GEN_237; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_239 = 8'hef == io_data_in[15:8] ? 8'hdf : _GEN_238; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_240 = 8'hf0 == io_data_in[15:8] ? 8'h8c : _GEN_239; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_241 = 8'hf1 == io_data_in[15:8] ? 8'ha1 : _GEN_240; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_242 = 8'hf2 == io_data_in[15:8] ? 8'h89 : _GEN_241; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_243 = 8'hf3 == io_data_in[15:8] ? 8'hd : _GEN_242; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_244 = 8'hf4 == io_data_in[15:8] ? 8'hbf : _GEN_243; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_245 = 8'hf5 == io_data_in[15:8] ? 8'he6 : _GEN_244; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_246 = 8'hf6 == io_data_in[15:8] ? 8'h42 : _GEN_245; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_247 = 8'hf7 == io_data_in[15:8] ? 8'h68 : _GEN_246; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_248 = 8'hf8 == io_data_in[15:8] ? 8'h41 : _GEN_247; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_249 = 8'hf9 == io_data_in[15:8] ? 8'h99 : _GEN_248; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_250 = 8'hfa == io_data_in[15:8] ? 8'h2d : _GEN_249; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_251 = 8'hfb == io_data_in[15:8] ? 8'hf : _GEN_250; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_252 = 8'hfc == io_data_in[15:8] ? 8'hb0 : _GEN_251; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_253 = 8'hfd == io_data_in[15:8] ? 8'h54 : _GEN_252; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_254 = 8'hfe == io_data_in[15:8] ? 8'hbb : _GEN_253; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  wire [7:0] _GEN_257 = 8'h1 == io_data_in[23:16] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_258 = 8'h2 == io_data_in[23:16] ? 8'h77 : _GEN_257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_259 = 8'h3 == io_data_in[23:16] ? 8'h7b : _GEN_258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_260 = 8'h4 == io_data_in[23:16] ? 8'hf2 : _GEN_259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_261 = 8'h5 == io_data_in[23:16] ? 8'h6b : _GEN_260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_262 = 8'h6 == io_data_in[23:16] ? 8'h6f : _GEN_261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_263 = 8'h7 == io_data_in[23:16] ? 8'hc5 : _GEN_262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_264 = 8'h8 == io_data_in[23:16] ? 8'h30 : _GEN_263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_265 = 8'h9 == io_data_in[23:16] ? 8'h1 : _GEN_264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_266 = 8'ha == io_data_in[23:16] ? 8'h67 : _GEN_265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_267 = 8'hb == io_data_in[23:16] ? 8'h2b : _GEN_266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_268 = 8'hc == io_data_in[23:16] ? 8'hfe : _GEN_267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_269 = 8'hd == io_data_in[23:16] ? 8'hd7 : _GEN_268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_270 = 8'he == io_data_in[23:16] ? 8'hab : _GEN_269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_271 = 8'hf == io_data_in[23:16] ? 8'h76 : _GEN_270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_272 = 8'h10 == io_data_in[23:16] ? 8'hca : _GEN_271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_273 = 8'h11 == io_data_in[23:16] ? 8'h82 : _GEN_272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_274 = 8'h12 == io_data_in[23:16] ? 8'hc9 : _GEN_273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_275 = 8'h13 == io_data_in[23:16] ? 8'h7d : _GEN_274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_276 = 8'h14 == io_data_in[23:16] ? 8'hfa : _GEN_275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_277 = 8'h15 == io_data_in[23:16] ? 8'h59 : _GEN_276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_278 = 8'h16 == io_data_in[23:16] ? 8'h47 : _GEN_277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_279 = 8'h17 == io_data_in[23:16] ? 8'hf0 : _GEN_278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_280 = 8'h18 == io_data_in[23:16] ? 8'had : _GEN_279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_281 = 8'h19 == io_data_in[23:16] ? 8'hd4 : _GEN_280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_282 = 8'h1a == io_data_in[23:16] ? 8'ha2 : _GEN_281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_283 = 8'h1b == io_data_in[23:16] ? 8'haf : _GEN_282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_284 = 8'h1c == io_data_in[23:16] ? 8'h9c : _GEN_283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_285 = 8'h1d == io_data_in[23:16] ? 8'ha4 : _GEN_284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_286 = 8'h1e == io_data_in[23:16] ? 8'h72 : _GEN_285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_287 = 8'h1f == io_data_in[23:16] ? 8'hc0 : _GEN_286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_288 = 8'h20 == io_data_in[23:16] ? 8'hb7 : _GEN_287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_289 = 8'h21 == io_data_in[23:16] ? 8'hfd : _GEN_288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_290 = 8'h22 == io_data_in[23:16] ? 8'h93 : _GEN_289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_291 = 8'h23 == io_data_in[23:16] ? 8'h26 : _GEN_290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_292 = 8'h24 == io_data_in[23:16] ? 8'h36 : _GEN_291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_293 = 8'h25 == io_data_in[23:16] ? 8'h3f : _GEN_292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_294 = 8'h26 == io_data_in[23:16] ? 8'hf7 : _GEN_293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_295 = 8'h27 == io_data_in[23:16] ? 8'hcc : _GEN_294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_296 = 8'h28 == io_data_in[23:16] ? 8'h34 : _GEN_295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_297 = 8'h29 == io_data_in[23:16] ? 8'ha5 : _GEN_296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_298 = 8'h2a == io_data_in[23:16] ? 8'he5 : _GEN_297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_299 = 8'h2b == io_data_in[23:16] ? 8'hf1 : _GEN_298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_300 = 8'h2c == io_data_in[23:16] ? 8'h71 : _GEN_299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_301 = 8'h2d == io_data_in[23:16] ? 8'hd8 : _GEN_300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_302 = 8'h2e == io_data_in[23:16] ? 8'h31 : _GEN_301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_303 = 8'h2f == io_data_in[23:16] ? 8'h15 : _GEN_302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_304 = 8'h30 == io_data_in[23:16] ? 8'h4 : _GEN_303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_305 = 8'h31 == io_data_in[23:16] ? 8'hc7 : _GEN_304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_306 = 8'h32 == io_data_in[23:16] ? 8'h23 : _GEN_305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_307 = 8'h33 == io_data_in[23:16] ? 8'hc3 : _GEN_306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_308 = 8'h34 == io_data_in[23:16] ? 8'h18 : _GEN_307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_309 = 8'h35 == io_data_in[23:16] ? 8'h96 : _GEN_308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_310 = 8'h36 == io_data_in[23:16] ? 8'h5 : _GEN_309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_311 = 8'h37 == io_data_in[23:16] ? 8'h9a : _GEN_310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_312 = 8'h38 == io_data_in[23:16] ? 8'h7 : _GEN_311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_313 = 8'h39 == io_data_in[23:16] ? 8'h12 : _GEN_312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_314 = 8'h3a == io_data_in[23:16] ? 8'h80 : _GEN_313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_315 = 8'h3b == io_data_in[23:16] ? 8'he2 : _GEN_314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_316 = 8'h3c == io_data_in[23:16] ? 8'heb : _GEN_315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_317 = 8'h3d == io_data_in[23:16] ? 8'h27 : _GEN_316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_318 = 8'h3e == io_data_in[23:16] ? 8'hb2 : _GEN_317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_319 = 8'h3f == io_data_in[23:16] ? 8'h75 : _GEN_318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_320 = 8'h40 == io_data_in[23:16] ? 8'h9 : _GEN_319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_321 = 8'h41 == io_data_in[23:16] ? 8'h83 : _GEN_320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_322 = 8'h42 == io_data_in[23:16] ? 8'h2c : _GEN_321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_323 = 8'h43 == io_data_in[23:16] ? 8'h1a : _GEN_322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_324 = 8'h44 == io_data_in[23:16] ? 8'h1b : _GEN_323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_325 = 8'h45 == io_data_in[23:16] ? 8'h6e : _GEN_324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_326 = 8'h46 == io_data_in[23:16] ? 8'h5a : _GEN_325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_327 = 8'h47 == io_data_in[23:16] ? 8'ha0 : _GEN_326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_328 = 8'h48 == io_data_in[23:16] ? 8'h52 : _GEN_327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_329 = 8'h49 == io_data_in[23:16] ? 8'h3b : _GEN_328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_330 = 8'h4a == io_data_in[23:16] ? 8'hd6 : _GEN_329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_331 = 8'h4b == io_data_in[23:16] ? 8'hb3 : _GEN_330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_332 = 8'h4c == io_data_in[23:16] ? 8'h29 : _GEN_331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_333 = 8'h4d == io_data_in[23:16] ? 8'he3 : _GEN_332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_334 = 8'h4e == io_data_in[23:16] ? 8'h2f : _GEN_333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_335 = 8'h4f == io_data_in[23:16] ? 8'h84 : _GEN_334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_336 = 8'h50 == io_data_in[23:16] ? 8'h53 : _GEN_335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_337 = 8'h51 == io_data_in[23:16] ? 8'hd1 : _GEN_336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_338 = 8'h52 == io_data_in[23:16] ? 8'h0 : _GEN_337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_339 = 8'h53 == io_data_in[23:16] ? 8'hed : _GEN_338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_340 = 8'h54 == io_data_in[23:16] ? 8'h20 : _GEN_339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_341 = 8'h55 == io_data_in[23:16] ? 8'hfc : _GEN_340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_342 = 8'h56 == io_data_in[23:16] ? 8'hb1 : _GEN_341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_343 = 8'h57 == io_data_in[23:16] ? 8'h5b : _GEN_342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_344 = 8'h58 == io_data_in[23:16] ? 8'h6a : _GEN_343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_345 = 8'h59 == io_data_in[23:16] ? 8'hcb : _GEN_344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_346 = 8'h5a == io_data_in[23:16] ? 8'hbe : _GEN_345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_347 = 8'h5b == io_data_in[23:16] ? 8'h39 : _GEN_346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_348 = 8'h5c == io_data_in[23:16] ? 8'h4a : _GEN_347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_349 = 8'h5d == io_data_in[23:16] ? 8'h4c : _GEN_348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_350 = 8'h5e == io_data_in[23:16] ? 8'h58 : _GEN_349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_351 = 8'h5f == io_data_in[23:16] ? 8'hcf : _GEN_350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_352 = 8'h60 == io_data_in[23:16] ? 8'hd0 : _GEN_351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_353 = 8'h61 == io_data_in[23:16] ? 8'hef : _GEN_352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_354 = 8'h62 == io_data_in[23:16] ? 8'haa : _GEN_353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_355 = 8'h63 == io_data_in[23:16] ? 8'hfb : _GEN_354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_356 = 8'h64 == io_data_in[23:16] ? 8'h43 : _GEN_355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_357 = 8'h65 == io_data_in[23:16] ? 8'h4d : _GEN_356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_358 = 8'h66 == io_data_in[23:16] ? 8'h33 : _GEN_357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_359 = 8'h67 == io_data_in[23:16] ? 8'h85 : _GEN_358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_360 = 8'h68 == io_data_in[23:16] ? 8'h45 : _GEN_359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_361 = 8'h69 == io_data_in[23:16] ? 8'hf9 : _GEN_360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_362 = 8'h6a == io_data_in[23:16] ? 8'h2 : _GEN_361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_363 = 8'h6b == io_data_in[23:16] ? 8'h7f : _GEN_362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_364 = 8'h6c == io_data_in[23:16] ? 8'h50 : _GEN_363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_365 = 8'h6d == io_data_in[23:16] ? 8'h3c : _GEN_364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_366 = 8'h6e == io_data_in[23:16] ? 8'h9f : _GEN_365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_367 = 8'h6f == io_data_in[23:16] ? 8'ha8 : _GEN_366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_368 = 8'h70 == io_data_in[23:16] ? 8'h51 : _GEN_367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_369 = 8'h71 == io_data_in[23:16] ? 8'ha3 : _GEN_368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_370 = 8'h72 == io_data_in[23:16] ? 8'h40 : _GEN_369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_371 = 8'h73 == io_data_in[23:16] ? 8'h8f : _GEN_370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_372 = 8'h74 == io_data_in[23:16] ? 8'h92 : _GEN_371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_373 = 8'h75 == io_data_in[23:16] ? 8'h9d : _GEN_372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_374 = 8'h76 == io_data_in[23:16] ? 8'h38 : _GEN_373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_375 = 8'h77 == io_data_in[23:16] ? 8'hf5 : _GEN_374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_376 = 8'h78 == io_data_in[23:16] ? 8'hbc : _GEN_375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_377 = 8'h79 == io_data_in[23:16] ? 8'hb6 : _GEN_376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_378 = 8'h7a == io_data_in[23:16] ? 8'hda : _GEN_377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_379 = 8'h7b == io_data_in[23:16] ? 8'h21 : _GEN_378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_380 = 8'h7c == io_data_in[23:16] ? 8'h10 : _GEN_379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_381 = 8'h7d == io_data_in[23:16] ? 8'hff : _GEN_380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_382 = 8'h7e == io_data_in[23:16] ? 8'hf3 : _GEN_381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_383 = 8'h7f == io_data_in[23:16] ? 8'hd2 : _GEN_382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_384 = 8'h80 == io_data_in[23:16] ? 8'hcd : _GEN_383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_385 = 8'h81 == io_data_in[23:16] ? 8'hc : _GEN_384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_386 = 8'h82 == io_data_in[23:16] ? 8'h13 : _GEN_385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_387 = 8'h83 == io_data_in[23:16] ? 8'hec : _GEN_386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_388 = 8'h84 == io_data_in[23:16] ? 8'h5f : _GEN_387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_389 = 8'h85 == io_data_in[23:16] ? 8'h97 : _GEN_388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_390 = 8'h86 == io_data_in[23:16] ? 8'h44 : _GEN_389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_391 = 8'h87 == io_data_in[23:16] ? 8'h17 : _GEN_390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_392 = 8'h88 == io_data_in[23:16] ? 8'hc4 : _GEN_391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_393 = 8'h89 == io_data_in[23:16] ? 8'ha7 : _GEN_392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_394 = 8'h8a == io_data_in[23:16] ? 8'h7e : _GEN_393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_395 = 8'h8b == io_data_in[23:16] ? 8'h3d : _GEN_394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_396 = 8'h8c == io_data_in[23:16] ? 8'h64 : _GEN_395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_397 = 8'h8d == io_data_in[23:16] ? 8'h5d : _GEN_396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_398 = 8'h8e == io_data_in[23:16] ? 8'h19 : _GEN_397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_399 = 8'h8f == io_data_in[23:16] ? 8'h73 : _GEN_398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_400 = 8'h90 == io_data_in[23:16] ? 8'h60 : _GEN_399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_401 = 8'h91 == io_data_in[23:16] ? 8'h81 : _GEN_400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_402 = 8'h92 == io_data_in[23:16] ? 8'h4f : _GEN_401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_403 = 8'h93 == io_data_in[23:16] ? 8'hdc : _GEN_402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_404 = 8'h94 == io_data_in[23:16] ? 8'h22 : _GEN_403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_405 = 8'h95 == io_data_in[23:16] ? 8'h2a : _GEN_404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_406 = 8'h96 == io_data_in[23:16] ? 8'h90 : _GEN_405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_407 = 8'h97 == io_data_in[23:16] ? 8'h88 : _GEN_406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_408 = 8'h98 == io_data_in[23:16] ? 8'h46 : _GEN_407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_409 = 8'h99 == io_data_in[23:16] ? 8'hee : _GEN_408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_410 = 8'h9a == io_data_in[23:16] ? 8'hb8 : _GEN_409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_411 = 8'h9b == io_data_in[23:16] ? 8'h14 : _GEN_410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_412 = 8'h9c == io_data_in[23:16] ? 8'hde : _GEN_411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_413 = 8'h9d == io_data_in[23:16] ? 8'h5e : _GEN_412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_414 = 8'h9e == io_data_in[23:16] ? 8'hb : _GEN_413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_415 = 8'h9f == io_data_in[23:16] ? 8'hdb : _GEN_414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_416 = 8'ha0 == io_data_in[23:16] ? 8'he0 : _GEN_415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_417 = 8'ha1 == io_data_in[23:16] ? 8'h32 : _GEN_416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_418 = 8'ha2 == io_data_in[23:16] ? 8'h3a : _GEN_417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_419 = 8'ha3 == io_data_in[23:16] ? 8'ha : _GEN_418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_420 = 8'ha4 == io_data_in[23:16] ? 8'h49 : _GEN_419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_421 = 8'ha5 == io_data_in[23:16] ? 8'h6 : _GEN_420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_422 = 8'ha6 == io_data_in[23:16] ? 8'h24 : _GEN_421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_423 = 8'ha7 == io_data_in[23:16] ? 8'h5c : _GEN_422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_424 = 8'ha8 == io_data_in[23:16] ? 8'hc2 : _GEN_423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_425 = 8'ha9 == io_data_in[23:16] ? 8'hd3 : _GEN_424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_426 = 8'haa == io_data_in[23:16] ? 8'hac : _GEN_425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_427 = 8'hab == io_data_in[23:16] ? 8'h62 : _GEN_426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_428 = 8'hac == io_data_in[23:16] ? 8'h91 : _GEN_427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_429 = 8'had == io_data_in[23:16] ? 8'h95 : _GEN_428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_430 = 8'hae == io_data_in[23:16] ? 8'he4 : _GEN_429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_431 = 8'haf == io_data_in[23:16] ? 8'h79 : _GEN_430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_432 = 8'hb0 == io_data_in[23:16] ? 8'he7 : _GEN_431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_433 = 8'hb1 == io_data_in[23:16] ? 8'hc8 : _GEN_432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_434 = 8'hb2 == io_data_in[23:16] ? 8'h37 : _GEN_433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_435 = 8'hb3 == io_data_in[23:16] ? 8'h6d : _GEN_434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_436 = 8'hb4 == io_data_in[23:16] ? 8'h8d : _GEN_435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_437 = 8'hb5 == io_data_in[23:16] ? 8'hd5 : _GEN_436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_438 = 8'hb6 == io_data_in[23:16] ? 8'h4e : _GEN_437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_439 = 8'hb7 == io_data_in[23:16] ? 8'ha9 : _GEN_438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_440 = 8'hb8 == io_data_in[23:16] ? 8'h6c : _GEN_439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_441 = 8'hb9 == io_data_in[23:16] ? 8'h56 : _GEN_440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_442 = 8'hba == io_data_in[23:16] ? 8'hf4 : _GEN_441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_443 = 8'hbb == io_data_in[23:16] ? 8'hea : _GEN_442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_444 = 8'hbc == io_data_in[23:16] ? 8'h65 : _GEN_443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_445 = 8'hbd == io_data_in[23:16] ? 8'h7a : _GEN_444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_446 = 8'hbe == io_data_in[23:16] ? 8'hae : _GEN_445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_447 = 8'hbf == io_data_in[23:16] ? 8'h8 : _GEN_446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_448 = 8'hc0 == io_data_in[23:16] ? 8'hba : _GEN_447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_449 = 8'hc1 == io_data_in[23:16] ? 8'h78 : _GEN_448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_450 = 8'hc2 == io_data_in[23:16] ? 8'h25 : _GEN_449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_451 = 8'hc3 == io_data_in[23:16] ? 8'h2e : _GEN_450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_452 = 8'hc4 == io_data_in[23:16] ? 8'h1c : _GEN_451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_453 = 8'hc5 == io_data_in[23:16] ? 8'ha6 : _GEN_452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_454 = 8'hc6 == io_data_in[23:16] ? 8'hb4 : _GEN_453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_455 = 8'hc7 == io_data_in[23:16] ? 8'hc6 : _GEN_454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_456 = 8'hc8 == io_data_in[23:16] ? 8'he8 : _GEN_455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_457 = 8'hc9 == io_data_in[23:16] ? 8'hdd : _GEN_456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_458 = 8'hca == io_data_in[23:16] ? 8'h74 : _GEN_457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_459 = 8'hcb == io_data_in[23:16] ? 8'h1f : _GEN_458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_460 = 8'hcc == io_data_in[23:16] ? 8'h4b : _GEN_459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_461 = 8'hcd == io_data_in[23:16] ? 8'hbd : _GEN_460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_462 = 8'hce == io_data_in[23:16] ? 8'h8b : _GEN_461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_463 = 8'hcf == io_data_in[23:16] ? 8'h8a : _GEN_462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_464 = 8'hd0 == io_data_in[23:16] ? 8'h70 : _GEN_463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_465 = 8'hd1 == io_data_in[23:16] ? 8'h3e : _GEN_464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_466 = 8'hd2 == io_data_in[23:16] ? 8'hb5 : _GEN_465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_467 = 8'hd3 == io_data_in[23:16] ? 8'h66 : _GEN_466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_468 = 8'hd4 == io_data_in[23:16] ? 8'h48 : _GEN_467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_469 = 8'hd5 == io_data_in[23:16] ? 8'h3 : _GEN_468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_470 = 8'hd6 == io_data_in[23:16] ? 8'hf6 : _GEN_469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_471 = 8'hd7 == io_data_in[23:16] ? 8'he : _GEN_470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_472 = 8'hd8 == io_data_in[23:16] ? 8'h61 : _GEN_471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_473 = 8'hd9 == io_data_in[23:16] ? 8'h35 : _GEN_472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_474 = 8'hda == io_data_in[23:16] ? 8'h57 : _GEN_473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_475 = 8'hdb == io_data_in[23:16] ? 8'hb9 : _GEN_474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_476 = 8'hdc == io_data_in[23:16] ? 8'h86 : _GEN_475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_477 = 8'hdd == io_data_in[23:16] ? 8'hc1 : _GEN_476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_478 = 8'hde == io_data_in[23:16] ? 8'h1d : _GEN_477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_479 = 8'hdf == io_data_in[23:16] ? 8'h9e : _GEN_478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_480 = 8'he0 == io_data_in[23:16] ? 8'he1 : _GEN_479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_481 = 8'he1 == io_data_in[23:16] ? 8'hf8 : _GEN_480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_482 = 8'he2 == io_data_in[23:16] ? 8'h98 : _GEN_481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_483 = 8'he3 == io_data_in[23:16] ? 8'h11 : _GEN_482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_484 = 8'he4 == io_data_in[23:16] ? 8'h69 : _GEN_483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_485 = 8'he5 == io_data_in[23:16] ? 8'hd9 : _GEN_484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_486 = 8'he6 == io_data_in[23:16] ? 8'h8e : _GEN_485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_487 = 8'he7 == io_data_in[23:16] ? 8'h94 : _GEN_486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_488 = 8'he8 == io_data_in[23:16] ? 8'h9b : _GEN_487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_489 = 8'he9 == io_data_in[23:16] ? 8'h1e : _GEN_488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_490 = 8'hea == io_data_in[23:16] ? 8'h87 : _GEN_489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_491 = 8'heb == io_data_in[23:16] ? 8'he9 : _GEN_490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_492 = 8'hec == io_data_in[23:16] ? 8'hce : _GEN_491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_493 = 8'hed == io_data_in[23:16] ? 8'h55 : _GEN_492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_494 = 8'hee == io_data_in[23:16] ? 8'h28 : _GEN_493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_495 = 8'hef == io_data_in[23:16] ? 8'hdf : _GEN_494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_496 = 8'hf0 == io_data_in[23:16] ? 8'h8c : _GEN_495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_497 = 8'hf1 == io_data_in[23:16] ? 8'ha1 : _GEN_496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_498 = 8'hf2 == io_data_in[23:16] ? 8'h89 : _GEN_497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_499 = 8'hf3 == io_data_in[23:16] ? 8'hd : _GEN_498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_500 = 8'hf4 == io_data_in[23:16] ? 8'hbf : _GEN_499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_501 = 8'hf5 == io_data_in[23:16] ? 8'he6 : _GEN_500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_502 = 8'hf6 == io_data_in[23:16] ? 8'h42 : _GEN_501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_503 = 8'hf7 == io_data_in[23:16] ? 8'h68 : _GEN_502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_504 = 8'hf8 == io_data_in[23:16] ? 8'h41 : _GEN_503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_505 = 8'hf9 == io_data_in[23:16] ? 8'h99 : _GEN_504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_506 = 8'hfa == io_data_in[23:16] ? 8'h2d : _GEN_505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_507 = 8'hfb == io_data_in[23:16] ? 8'hf : _GEN_506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_508 = 8'hfc == io_data_in[23:16] ? 8'hb0 : _GEN_507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_509 = 8'hfd == io_data_in[23:16] ? 8'h54 : _GEN_508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_510 = 8'hfe == io_data_in[23:16] ? 8'hbb : _GEN_509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_511 = 8'hff == io_data_in[23:16] ? 8'h16 : _GEN_510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [15:0] io_data_out_lo = {_GEN_511,io_data_out_a_io_data_out}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_513 = 8'h1 == io_data_in[7:0] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_514 = 8'h2 == io_data_in[7:0] ? 8'h77 : _GEN_513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_515 = 8'h3 == io_data_in[7:0] ? 8'h7b : _GEN_514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_516 = 8'h4 == io_data_in[7:0] ? 8'hf2 : _GEN_515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_517 = 8'h5 == io_data_in[7:0] ? 8'h6b : _GEN_516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_518 = 8'h6 == io_data_in[7:0] ? 8'h6f : _GEN_517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_519 = 8'h7 == io_data_in[7:0] ? 8'hc5 : _GEN_518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_520 = 8'h8 == io_data_in[7:0] ? 8'h30 : _GEN_519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_521 = 8'h9 == io_data_in[7:0] ? 8'h1 : _GEN_520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_522 = 8'ha == io_data_in[7:0] ? 8'h67 : _GEN_521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_523 = 8'hb == io_data_in[7:0] ? 8'h2b : _GEN_522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_524 = 8'hc == io_data_in[7:0] ? 8'hfe : _GEN_523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_525 = 8'hd == io_data_in[7:0] ? 8'hd7 : _GEN_524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_526 = 8'he == io_data_in[7:0] ? 8'hab : _GEN_525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_527 = 8'hf == io_data_in[7:0] ? 8'h76 : _GEN_526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_528 = 8'h10 == io_data_in[7:0] ? 8'hca : _GEN_527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_529 = 8'h11 == io_data_in[7:0] ? 8'h82 : _GEN_528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_530 = 8'h12 == io_data_in[7:0] ? 8'hc9 : _GEN_529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_531 = 8'h13 == io_data_in[7:0] ? 8'h7d : _GEN_530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_532 = 8'h14 == io_data_in[7:0] ? 8'hfa : _GEN_531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_533 = 8'h15 == io_data_in[7:0] ? 8'h59 : _GEN_532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_534 = 8'h16 == io_data_in[7:0] ? 8'h47 : _GEN_533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_535 = 8'h17 == io_data_in[7:0] ? 8'hf0 : _GEN_534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_536 = 8'h18 == io_data_in[7:0] ? 8'had : _GEN_535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_537 = 8'h19 == io_data_in[7:0] ? 8'hd4 : _GEN_536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_538 = 8'h1a == io_data_in[7:0] ? 8'ha2 : _GEN_537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_539 = 8'h1b == io_data_in[7:0] ? 8'haf : _GEN_538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_540 = 8'h1c == io_data_in[7:0] ? 8'h9c : _GEN_539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_541 = 8'h1d == io_data_in[7:0] ? 8'ha4 : _GEN_540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_542 = 8'h1e == io_data_in[7:0] ? 8'h72 : _GEN_541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_543 = 8'h1f == io_data_in[7:0] ? 8'hc0 : _GEN_542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_544 = 8'h20 == io_data_in[7:0] ? 8'hb7 : _GEN_543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_545 = 8'h21 == io_data_in[7:0] ? 8'hfd : _GEN_544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_546 = 8'h22 == io_data_in[7:0] ? 8'h93 : _GEN_545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_547 = 8'h23 == io_data_in[7:0] ? 8'h26 : _GEN_546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_548 = 8'h24 == io_data_in[7:0] ? 8'h36 : _GEN_547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_549 = 8'h25 == io_data_in[7:0] ? 8'h3f : _GEN_548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_550 = 8'h26 == io_data_in[7:0] ? 8'hf7 : _GEN_549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_551 = 8'h27 == io_data_in[7:0] ? 8'hcc : _GEN_550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_552 = 8'h28 == io_data_in[7:0] ? 8'h34 : _GEN_551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_553 = 8'h29 == io_data_in[7:0] ? 8'ha5 : _GEN_552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_554 = 8'h2a == io_data_in[7:0] ? 8'he5 : _GEN_553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_555 = 8'h2b == io_data_in[7:0] ? 8'hf1 : _GEN_554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_556 = 8'h2c == io_data_in[7:0] ? 8'h71 : _GEN_555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_557 = 8'h2d == io_data_in[7:0] ? 8'hd8 : _GEN_556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_558 = 8'h2e == io_data_in[7:0] ? 8'h31 : _GEN_557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_559 = 8'h2f == io_data_in[7:0] ? 8'h15 : _GEN_558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_560 = 8'h30 == io_data_in[7:0] ? 8'h4 : _GEN_559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_561 = 8'h31 == io_data_in[7:0] ? 8'hc7 : _GEN_560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_562 = 8'h32 == io_data_in[7:0] ? 8'h23 : _GEN_561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_563 = 8'h33 == io_data_in[7:0] ? 8'hc3 : _GEN_562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_564 = 8'h34 == io_data_in[7:0] ? 8'h18 : _GEN_563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_565 = 8'h35 == io_data_in[7:0] ? 8'h96 : _GEN_564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_566 = 8'h36 == io_data_in[7:0] ? 8'h5 : _GEN_565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_567 = 8'h37 == io_data_in[7:0] ? 8'h9a : _GEN_566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_568 = 8'h38 == io_data_in[7:0] ? 8'h7 : _GEN_567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_569 = 8'h39 == io_data_in[7:0] ? 8'h12 : _GEN_568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_570 = 8'h3a == io_data_in[7:0] ? 8'h80 : _GEN_569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_571 = 8'h3b == io_data_in[7:0] ? 8'he2 : _GEN_570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_572 = 8'h3c == io_data_in[7:0] ? 8'heb : _GEN_571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_573 = 8'h3d == io_data_in[7:0] ? 8'h27 : _GEN_572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_574 = 8'h3e == io_data_in[7:0] ? 8'hb2 : _GEN_573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_575 = 8'h3f == io_data_in[7:0] ? 8'h75 : _GEN_574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_576 = 8'h40 == io_data_in[7:0] ? 8'h9 : _GEN_575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_577 = 8'h41 == io_data_in[7:0] ? 8'h83 : _GEN_576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_578 = 8'h42 == io_data_in[7:0] ? 8'h2c : _GEN_577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_579 = 8'h43 == io_data_in[7:0] ? 8'h1a : _GEN_578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_580 = 8'h44 == io_data_in[7:0] ? 8'h1b : _GEN_579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_581 = 8'h45 == io_data_in[7:0] ? 8'h6e : _GEN_580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_582 = 8'h46 == io_data_in[7:0] ? 8'h5a : _GEN_581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_583 = 8'h47 == io_data_in[7:0] ? 8'ha0 : _GEN_582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_584 = 8'h48 == io_data_in[7:0] ? 8'h52 : _GEN_583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_585 = 8'h49 == io_data_in[7:0] ? 8'h3b : _GEN_584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_586 = 8'h4a == io_data_in[7:0] ? 8'hd6 : _GEN_585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_587 = 8'h4b == io_data_in[7:0] ? 8'hb3 : _GEN_586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_588 = 8'h4c == io_data_in[7:0] ? 8'h29 : _GEN_587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_589 = 8'h4d == io_data_in[7:0] ? 8'he3 : _GEN_588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_590 = 8'h4e == io_data_in[7:0] ? 8'h2f : _GEN_589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_591 = 8'h4f == io_data_in[7:0] ? 8'h84 : _GEN_590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_592 = 8'h50 == io_data_in[7:0] ? 8'h53 : _GEN_591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_593 = 8'h51 == io_data_in[7:0] ? 8'hd1 : _GEN_592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_594 = 8'h52 == io_data_in[7:0] ? 8'h0 : _GEN_593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_595 = 8'h53 == io_data_in[7:0] ? 8'hed : _GEN_594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_596 = 8'h54 == io_data_in[7:0] ? 8'h20 : _GEN_595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_597 = 8'h55 == io_data_in[7:0] ? 8'hfc : _GEN_596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_598 = 8'h56 == io_data_in[7:0] ? 8'hb1 : _GEN_597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_599 = 8'h57 == io_data_in[7:0] ? 8'h5b : _GEN_598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_600 = 8'h58 == io_data_in[7:0] ? 8'h6a : _GEN_599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_601 = 8'h59 == io_data_in[7:0] ? 8'hcb : _GEN_600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_602 = 8'h5a == io_data_in[7:0] ? 8'hbe : _GEN_601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_603 = 8'h5b == io_data_in[7:0] ? 8'h39 : _GEN_602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_604 = 8'h5c == io_data_in[7:0] ? 8'h4a : _GEN_603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_605 = 8'h5d == io_data_in[7:0] ? 8'h4c : _GEN_604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_606 = 8'h5e == io_data_in[7:0] ? 8'h58 : _GEN_605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_607 = 8'h5f == io_data_in[7:0] ? 8'hcf : _GEN_606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_608 = 8'h60 == io_data_in[7:0] ? 8'hd0 : _GEN_607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_609 = 8'h61 == io_data_in[7:0] ? 8'hef : _GEN_608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_610 = 8'h62 == io_data_in[7:0] ? 8'haa : _GEN_609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_611 = 8'h63 == io_data_in[7:0] ? 8'hfb : _GEN_610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_612 = 8'h64 == io_data_in[7:0] ? 8'h43 : _GEN_611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_613 = 8'h65 == io_data_in[7:0] ? 8'h4d : _GEN_612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_614 = 8'h66 == io_data_in[7:0] ? 8'h33 : _GEN_613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_615 = 8'h67 == io_data_in[7:0] ? 8'h85 : _GEN_614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_616 = 8'h68 == io_data_in[7:0] ? 8'h45 : _GEN_615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_617 = 8'h69 == io_data_in[7:0] ? 8'hf9 : _GEN_616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_618 = 8'h6a == io_data_in[7:0] ? 8'h2 : _GEN_617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_619 = 8'h6b == io_data_in[7:0] ? 8'h7f : _GEN_618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_620 = 8'h6c == io_data_in[7:0] ? 8'h50 : _GEN_619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_621 = 8'h6d == io_data_in[7:0] ? 8'h3c : _GEN_620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_622 = 8'h6e == io_data_in[7:0] ? 8'h9f : _GEN_621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_623 = 8'h6f == io_data_in[7:0] ? 8'ha8 : _GEN_622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_624 = 8'h70 == io_data_in[7:0] ? 8'h51 : _GEN_623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_625 = 8'h71 == io_data_in[7:0] ? 8'ha3 : _GEN_624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_626 = 8'h72 == io_data_in[7:0] ? 8'h40 : _GEN_625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_627 = 8'h73 == io_data_in[7:0] ? 8'h8f : _GEN_626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_628 = 8'h74 == io_data_in[7:0] ? 8'h92 : _GEN_627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_629 = 8'h75 == io_data_in[7:0] ? 8'h9d : _GEN_628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_630 = 8'h76 == io_data_in[7:0] ? 8'h38 : _GEN_629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_631 = 8'h77 == io_data_in[7:0] ? 8'hf5 : _GEN_630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_632 = 8'h78 == io_data_in[7:0] ? 8'hbc : _GEN_631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_633 = 8'h79 == io_data_in[7:0] ? 8'hb6 : _GEN_632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_634 = 8'h7a == io_data_in[7:0] ? 8'hda : _GEN_633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_635 = 8'h7b == io_data_in[7:0] ? 8'h21 : _GEN_634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_636 = 8'h7c == io_data_in[7:0] ? 8'h10 : _GEN_635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_637 = 8'h7d == io_data_in[7:0] ? 8'hff : _GEN_636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_638 = 8'h7e == io_data_in[7:0] ? 8'hf3 : _GEN_637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_639 = 8'h7f == io_data_in[7:0] ? 8'hd2 : _GEN_638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_640 = 8'h80 == io_data_in[7:0] ? 8'hcd : _GEN_639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_641 = 8'h81 == io_data_in[7:0] ? 8'hc : _GEN_640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_642 = 8'h82 == io_data_in[7:0] ? 8'h13 : _GEN_641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_643 = 8'h83 == io_data_in[7:0] ? 8'hec : _GEN_642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_644 = 8'h84 == io_data_in[7:0] ? 8'h5f : _GEN_643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_645 = 8'h85 == io_data_in[7:0] ? 8'h97 : _GEN_644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_646 = 8'h86 == io_data_in[7:0] ? 8'h44 : _GEN_645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_647 = 8'h87 == io_data_in[7:0] ? 8'h17 : _GEN_646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_648 = 8'h88 == io_data_in[7:0] ? 8'hc4 : _GEN_647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_649 = 8'h89 == io_data_in[7:0] ? 8'ha7 : _GEN_648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_650 = 8'h8a == io_data_in[7:0] ? 8'h7e : _GEN_649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_651 = 8'h8b == io_data_in[7:0] ? 8'h3d : _GEN_650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_652 = 8'h8c == io_data_in[7:0] ? 8'h64 : _GEN_651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_653 = 8'h8d == io_data_in[7:0] ? 8'h5d : _GEN_652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_654 = 8'h8e == io_data_in[7:0] ? 8'h19 : _GEN_653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_655 = 8'h8f == io_data_in[7:0] ? 8'h73 : _GEN_654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_656 = 8'h90 == io_data_in[7:0] ? 8'h60 : _GEN_655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_657 = 8'h91 == io_data_in[7:0] ? 8'h81 : _GEN_656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_658 = 8'h92 == io_data_in[7:0] ? 8'h4f : _GEN_657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_659 = 8'h93 == io_data_in[7:0] ? 8'hdc : _GEN_658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_660 = 8'h94 == io_data_in[7:0] ? 8'h22 : _GEN_659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_661 = 8'h95 == io_data_in[7:0] ? 8'h2a : _GEN_660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_662 = 8'h96 == io_data_in[7:0] ? 8'h90 : _GEN_661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_663 = 8'h97 == io_data_in[7:0] ? 8'h88 : _GEN_662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_664 = 8'h98 == io_data_in[7:0] ? 8'h46 : _GEN_663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_665 = 8'h99 == io_data_in[7:0] ? 8'hee : _GEN_664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_666 = 8'h9a == io_data_in[7:0] ? 8'hb8 : _GEN_665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_667 = 8'h9b == io_data_in[7:0] ? 8'h14 : _GEN_666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_668 = 8'h9c == io_data_in[7:0] ? 8'hde : _GEN_667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_669 = 8'h9d == io_data_in[7:0] ? 8'h5e : _GEN_668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_670 = 8'h9e == io_data_in[7:0] ? 8'hb : _GEN_669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_671 = 8'h9f == io_data_in[7:0] ? 8'hdb : _GEN_670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_672 = 8'ha0 == io_data_in[7:0] ? 8'he0 : _GEN_671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_673 = 8'ha1 == io_data_in[7:0] ? 8'h32 : _GEN_672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_674 = 8'ha2 == io_data_in[7:0] ? 8'h3a : _GEN_673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_675 = 8'ha3 == io_data_in[7:0] ? 8'ha : _GEN_674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_676 = 8'ha4 == io_data_in[7:0] ? 8'h49 : _GEN_675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_677 = 8'ha5 == io_data_in[7:0] ? 8'h6 : _GEN_676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_678 = 8'ha6 == io_data_in[7:0] ? 8'h24 : _GEN_677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_679 = 8'ha7 == io_data_in[7:0] ? 8'h5c : _GEN_678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_680 = 8'ha8 == io_data_in[7:0] ? 8'hc2 : _GEN_679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_681 = 8'ha9 == io_data_in[7:0] ? 8'hd3 : _GEN_680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_682 = 8'haa == io_data_in[7:0] ? 8'hac : _GEN_681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_683 = 8'hab == io_data_in[7:0] ? 8'h62 : _GEN_682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_684 = 8'hac == io_data_in[7:0] ? 8'h91 : _GEN_683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_685 = 8'had == io_data_in[7:0] ? 8'h95 : _GEN_684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_686 = 8'hae == io_data_in[7:0] ? 8'he4 : _GEN_685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_687 = 8'haf == io_data_in[7:0] ? 8'h79 : _GEN_686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_688 = 8'hb0 == io_data_in[7:0] ? 8'he7 : _GEN_687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_689 = 8'hb1 == io_data_in[7:0] ? 8'hc8 : _GEN_688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_690 = 8'hb2 == io_data_in[7:0] ? 8'h37 : _GEN_689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_691 = 8'hb3 == io_data_in[7:0] ? 8'h6d : _GEN_690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_692 = 8'hb4 == io_data_in[7:0] ? 8'h8d : _GEN_691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_693 = 8'hb5 == io_data_in[7:0] ? 8'hd5 : _GEN_692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_694 = 8'hb6 == io_data_in[7:0] ? 8'h4e : _GEN_693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_695 = 8'hb7 == io_data_in[7:0] ? 8'ha9 : _GEN_694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_696 = 8'hb8 == io_data_in[7:0] ? 8'h6c : _GEN_695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_697 = 8'hb9 == io_data_in[7:0] ? 8'h56 : _GEN_696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_698 = 8'hba == io_data_in[7:0] ? 8'hf4 : _GEN_697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_699 = 8'hbb == io_data_in[7:0] ? 8'hea : _GEN_698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_700 = 8'hbc == io_data_in[7:0] ? 8'h65 : _GEN_699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_701 = 8'hbd == io_data_in[7:0] ? 8'h7a : _GEN_700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_702 = 8'hbe == io_data_in[7:0] ? 8'hae : _GEN_701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_703 = 8'hbf == io_data_in[7:0] ? 8'h8 : _GEN_702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_704 = 8'hc0 == io_data_in[7:0] ? 8'hba : _GEN_703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_705 = 8'hc1 == io_data_in[7:0] ? 8'h78 : _GEN_704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_706 = 8'hc2 == io_data_in[7:0] ? 8'h25 : _GEN_705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_707 = 8'hc3 == io_data_in[7:0] ? 8'h2e : _GEN_706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_708 = 8'hc4 == io_data_in[7:0] ? 8'h1c : _GEN_707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_709 = 8'hc5 == io_data_in[7:0] ? 8'ha6 : _GEN_708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_710 = 8'hc6 == io_data_in[7:0] ? 8'hb4 : _GEN_709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_711 = 8'hc7 == io_data_in[7:0] ? 8'hc6 : _GEN_710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_712 = 8'hc8 == io_data_in[7:0] ? 8'he8 : _GEN_711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_713 = 8'hc9 == io_data_in[7:0] ? 8'hdd : _GEN_712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_714 = 8'hca == io_data_in[7:0] ? 8'h74 : _GEN_713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_715 = 8'hcb == io_data_in[7:0] ? 8'h1f : _GEN_714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_716 = 8'hcc == io_data_in[7:0] ? 8'h4b : _GEN_715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_717 = 8'hcd == io_data_in[7:0] ? 8'hbd : _GEN_716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_718 = 8'hce == io_data_in[7:0] ? 8'h8b : _GEN_717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_719 = 8'hcf == io_data_in[7:0] ? 8'h8a : _GEN_718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_720 = 8'hd0 == io_data_in[7:0] ? 8'h70 : _GEN_719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_721 = 8'hd1 == io_data_in[7:0] ? 8'h3e : _GEN_720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_722 = 8'hd2 == io_data_in[7:0] ? 8'hb5 : _GEN_721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_723 = 8'hd3 == io_data_in[7:0] ? 8'h66 : _GEN_722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_724 = 8'hd4 == io_data_in[7:0] ? 8'h48 : _GEN_723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_725 = 8'hd5 == io_data_in[7:0] ? 8'h3 : _GEN_724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_726 = 8'hd6 == io_data_in[7:0] ? 8'hf6 : _GEN_725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_727 = 8'hd7 == io_data_in[7:0] ? 8'he : _GEN_726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_728 = 8'hd8 == io_data_in[7:0] ? 8'h61 : _GEN_727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_729 = 8'hd9 == io_data_in[7:0] ? 8'h35 : _GEN_728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_730 = 8'hda == io_data_in[7:0] ? 8'h57 : _GEN_729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_731 = 8'hdb == io_data_in[7:0] ? 8'hb9 : _GEN_730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_732 = 8'hdc == io_data_in[7:0] ? 8'h86 : _GEN_731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_733 = 8'hdd == io_data_in[7:0] ? 8'hc1 : _GEN_732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_734 = 8'hde == io_data_in[7:0] ? 8'h1d : _GEN_733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_735 = 8'hdf == io_data_in[7:0] ? 8'h9e : _GEN_734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_736 = 8'he0 == io_data_in[7:0] ? 8'he1 : _GEN_735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_737 = 8'he1 == io_data_in[7:0] ? 8'hf8 : _GEN_736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_738 = 8'he2 == io_data_in[7:0] ? 8'h98 : _GEN_737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_739 = 8'he3 == io_data_in[7:0] ? 8'h11 : _GEN_738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_740 = 8'he4 == io_data_in[7:0] ? 8'h69 : _GEN_739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_741 = 8'he5 == io_data_in[7:0] ? 8'hd9 : _GEN_740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_742 = 8'he6 == io_data_in[7:0] ? 8'h8e : _GEN_741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_743 = 8'he7 == io_data_in[7:0] ? 8'h94 : _GEN_742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_744 = 8'he8 == io_data_in[7:0] ? 8'h9b : _GEN_743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_745 = 8'he9 == io_data_in[7:0] ? 8'h1e : _GEN_744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_746 = 8'hea == io_data_in[7:0] ? 8'h87 : _GEN_745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_747 = 8'heb == io_data_in[7:0] ? 8'he9 : _GEN_746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_748 = 8'hec == io_data_in[7:0] ? 8'hce : _GEN_747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_749 = 8'hed == io_data_in[7:0] ? 8'h55 : _GEN_748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_750 = 8'hee == io_data_in[7:0] ? 8'h28 : _GEN_749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_751 = 8'hef == io_data_in[7:0] ? 8'hdf : _GEN_750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_752 = 8'hf0 == io_data_in[7:0] ? 8'h8c : _GEN_751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_753 = 8'hf1 == io_data_in[7:0] ? 8'ha1 : _GEN_752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_754 = 8'hf2 == io_data_in[7:0] ? 8'h89 : _GEN_753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_755 = 8'hf3 == io_data_in[7:0] ? 8'hd : _GEN_754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_756 = 8'hf4 == io_data_in[7:0] ? 8'hbf : _GEN_755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_757 = 8'hf5 == io_data_in[7:0] ? 8'he6 : _GEN_756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_758 = 8'hf6 == io_data_in[7:0] ? 8'h42 : _GEN_757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_759 = 8'hf7 == io_data_in[7:0] ? 8'h68 : _GEN_758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_760 = 8'hf8 == io_data_in[7:0] ? 8'h41 : _GEN_759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_761 = 8'hf9 == io_data_in[7:0] ? 8'h99 : _GEN_760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_762 = 8'hfa == io_data_in[7:0] ? 8'h2d : _GEN_761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_763 = 8'hfb == io_data_in[7:0] ? 8'hf : _GEN_762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_764 = 8'hfc == io_data_in[7:0] ? 8'hb0 : _GEN_763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_765 = 8'hfd == io_data_in[7:0] ? 8'h54 : _GEN_764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_766 = 8'hfe == io_data_in[7:0] ? 8'hbb : _GEN_765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_767 = 8'hff == io_data_in[7:0] ? 8'h16 : _GEN_766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_769 = 8'h1 == io_data_in[31:24] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_770 = 8'h2 == io_data_in[31:24] ? 8'h77 : _GEN_769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_771 = 8'h3 == io_data_in[31:24] ? 8'h7b : _GEN_770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_772 = 8'h4 == io_data_in[31:24] ? 8'hf2 : _GEN_771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_773 = 8'h5 == io_data_in[31:24] ? 8'h6b : _GEN_772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_774 = 8'h6 == io_data_in[31:24] ? 8'h6f : _GEN_773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_775 = 8'h7 == io_data_in[31:24] ? 8'hc5 : _GEN_774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_776 = 8'h8 == io_data_in[31:24] ? 8'h30 : _GEN_775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_777 = 8'h9 == io_data_in[31:24] ? 8'h1 : _GEN_776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_778 = 8'ha == io_data_in[31:24] ? 8'h67 : _GEN_777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_779 = 8'hb == io_data_in[31:24] ? 8'h2b : _GEN_778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_780 = 8'hc == io_data_in[31:24] ? 8'hfe : _GEN_779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_781 = 8'hd == io_data_in[31:24] ? 8'hd7 : _GEN_780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_782 = 8'he == io_data_in[31:24] ? 8'hab : _GEN_781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_783 = 8'hf == io_data_in[31:24] ? 8'h76 : _GEN_782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_784 = 8'h10 == io_data_in[31:24] ? 8'hca : _GEN_783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_785 = 8'h11 == io_data_in[31:24] ? 8'h82 : _GEN_784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_786 = 8'h12 == io_data_in[31:24] ? 8'hc9 : _GEN_785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_787 = 8'h13 == io_data_in[31:24] ? 8'h7d : _GEN_786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_788 = 8'h14 == io_data_in[31:24] ? 8'hfa : _GEN_787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_789 = 8'h15 == io_data_in[31:24] ? 8'h59 : _GEN_788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_790 = 8'h16 == io_data_in[31:24] ? 8'h47 : _GEN_789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_791 = 8'h17 == io_data_in[31:24] ? 8'hf0 : _GEN_790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_792 = 8'h18 == io_data_in[31:24] ? 8'had : _GEN_791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_793 = 8'h19 == io_data_in[31:24] ? 8'hd4 : _GEN_792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_794 = 8'h1a == io_data_in[31:24] ? 8'ha2 : _GEN_793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_795 = 8'h1b == io_data_in[31:24] ? 8'haf : _GEN_794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_796 = 8'h1c == io_data_in[31:24] ? 8'h9c : _GEN_795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_797 = 8'h1d == io_data_in[31:24] ? 8'ha4 : _GEN_796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_798 = 8'h1e == io_data_in[31:24] ? 8'h72 : _GEN_797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_799 = 8'h1f == io_data_in[31:24] ? 8'hc0 : _GEN_798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_800 = 8'h20 == io_data_in[31:24] ? 8'hb7 : _GEN_799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_801 = 8'h21 == io_data_in[31:24] ? 8'hfd : _GEN_800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_802 = 8'h22 == io_data_in[31:24] ? 8'h93 : _GEN_801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_803 = 8'h23 == io_data_in[31:24] ? 8'h26 : _GEN_802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_804 = 8'h24 == io_data_in[31:24] ? 8'h36 : _GEN_803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_805 = 8'h25 == io_data_in[31:24] ? 8'h3f : _GEN_804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_806 = 8'h26 == io_data_in[31:24] ? 8'hf7 : _GEN_805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_807 = 8'h27 == io_data_in[31:24] ? 8'hcc : _GEN_806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_808 = 8'h28 == io_data_in[31:24] ? 8'h34 : _GEN_807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_809 = 8'h29 == io_data_in[31:24] ? 8'ha5 : _GEN_808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_810 = 8'h2a == io_data_in[31:24] ? 8'he5 : _GEN_809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_811 = 8'h2b == io_data_in[31:24] ? 8'hf1 : _GEN_810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_812 = 8'h2c == io_data_in[31:24] ? 8'h71 : _GEN_811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_813 = 8'h2d == io_data_in[31:24] ? 8'hd8 : _GEN_812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_814 = 8'h2e == io_data_in[31:24] ? 8'h31 : _GEN_813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_815 = 8'h2f == io_data_in[31:24] ? 8'h15 : _GEN_814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_816 = 8'h30 == io_data_in[31:24] ? 8'h4 : _GEN_815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_817 = 8'h31 == io_data_in[31:24] ? 8'hc7 : _GEN_816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_818 = 8'h32 == io_data_in[31:24] ? 8'h23 : _GEN_817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_819 = 8'h33 == io_data_in[31:24] ? 8'hc3 : _GEN_818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_820 = 8'h34 == io_data_in[31:24] ? 8'h18 : _GEN_819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_821 = 8'h35 == io_data_in[31:24] ? 8'h96 : _GEN_820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_822 = 8'h36 == io_data_in[31:24] ? 8'h5 : _GEN_821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_823 = 8'h37 == io_data_in[31:24] ? 8'h9a : _GEN_822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_824 = 8'h38 == io_data_in[31:24] ? 8'h7 : _GEN_823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_825 = 8'h39 == io_data_in[31:24] ? 8'h12 : _GEN_824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_826 = 8'h3a == io_data_in[31:24] ? 8'h80 : _GEN_825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_827 = 8'h3b == io_data_in[31:24] ? 8'he2 : _GEN_826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_828 = 8'h3c == io_data_in[31:24] ? 8'heb : _GEN_827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_829 = 8'h3d == io_data_in[31:24] ? 8'h27 : _GEN_828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_830 = 8'h3e == io_data_in[31:24] ? 8'hb2 : _GEN_829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_831 = 8'h3f == io_data_in[31:24] ? 8'h75 : _GEN_830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_832 = 8'h40 == io_data_in[31:24] ? 8'h9 : _GEN_831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_833 = 8'h41 == io_data_in[31:24] ? 8'h83 : _GEN_832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_834 = 8'h42 == io_data_in[31:24] ? 8'h2c : _GEN_833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_835 = 8'h43 == io_data_in[31:24] ? 8'h1a : _GEN_834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_836 = 8'h44 == io_data_in[31:24] ? 8'h1b : _GEN_835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_837 = 8'h45 == io_data_in[31:24] ? 8'h6e : _GEN_836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_838 = 8'h46 == io_data_in[31:24] ? 8'h5a : _GEN_837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_839 = 8'h47 == io_data_in[31:24] ? 8'ha0 : _GEN_838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_840 = 8'h48 == io_data_in[31:24] ? 8'h52 : _GEN_839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_841 = 8'h49 == io_data_in[31:24] ? 8'h3b : _GEN_840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_842 = 8'h4a == io_data_in[31:24] ? 8'hd6 : _GEN_841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_843 = 8'h4b == io_data_in[31:24] ? 8'hb3 : _GEN_842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_844 = 8'h4c == io_data_in[31:24] ? 8'h29 : _GEN_843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_845 = 8'h4d == io_data_in[31:24] ? 8'he3 : _GEN_844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_846 = 8'h4e == io_data_in[31:24] ? 8'h2f : _GEN_845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_847 = 8'h4f == io_data_in[31:24] ? 8'h84 : _GEN_846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_848 = 8'h50 == io_data_in[31:24] ? 8'h53 : _GEN_847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_849 = 8'h51 == io_data_in[31:24] ? 8'hd1 : _GEN_848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_850 = 8'h52 == io_data_in[31:24] ? 8'h0 : _GEN_849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_851 = 8'h53 == io_data_in[31:24] ? 8'hed : _GEN_850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_852 = 8'h54 == io_data_in[31:24] ? 8'h20 : _GEN_851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_853 = 8'h55 == io_data_in[31:24] ? 8'hfc : _GEN_852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_854 = 8'h56 == io_data_in[31:24] ? 8'hb1 : _GEN_853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_855 = 8'h57 == io_data_in[31:24] ? 8'h5b : _GEN_854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_856 = 8'h58 == io_data_in[31:24] ? 8'h6a : _GEN_855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_857 = 8'h59 == io_data_in[31:24] ? 8'hcb : _GEN_856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_858 = 8'h5a == io_data_in[31:24] ? 8'hbe : _GEN_857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_859 = 8'h5b == io_data_in[31:24] ? 8'h39 : _GEN_858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_860 = 8'h5c == io_data_in[31:24] ? 8'h4a : _GEN_859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_861 = 8'h5d == io_data_in[31:24] ? 8'h4c : _GEN_860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_862 = 8'h5e == io_data_in[31:24] ? 8'h58 : _GEN_861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_863 = 8'h5f == io_data_in[31:24] ? 8'hcf : _GEN_862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_864 = 8'h60 == io_data_in[31:24] ? 8'hd0 : _GEN_863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_865 = 8'h61 == io_data_in[31:24] ? 8'hef : _GEN_864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_866 = 8'h62 == io_data_in[31:24] ? 8'haa : _GEN_865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_867 = 8'h63 == io_data_in[31:24] ? 8'hfb : _GEN_866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_868 = 8'h64 == io_data_in[31:24] ? 8'h43 : _GEN_867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_869 = 8'h65 == io_data_in[31:24] ? 8'h4d : _GEN_868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_870 = 8'h66 == io_data_in[31:24] ? 8'h33 : _GEN_869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_871 = 8'h67 == io_data_in[31:24] ? 8'h85 : _GEN_870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_872 = 8'h68 == io_data_in[31:24] ? 8'h45 : _GEN_871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_873 = 8'h69 == io_data_in[31:24] ? 8'hf9 : _GEN_872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_874 = 8'h6a == io_data_in[31:24] ? 8'h2 : _GEN_873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_875 = 8'h6b == io_data_in[31:24] ? 8'h7f : _GEN_874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_876 = 8'h6c == io_data_in[31:24] ? 8'h50 : _GEN_875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_877 = 8'h6d == io_data_in[31:24] ? 8'h3c : _GEN_876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_878 = 8'h6e == io_data_in[31:24] ? 8'h9f : _GEN_877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_879 = 8'h6f == io_data_in[31:24] ? 8'ha8 : _GEN_878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_880 = 8'h70 == io_data_in[31:24] ? 8'h51 : _GEN_879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_881 = 8'h71 == io_data_in[31:24] ? 8'ha3 : _GEN_880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_882 = 8'h72 == io_data_in[31:24] ? 8'h40 : _GEN_881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_883 = 8'h73 == io_data_in[31:24] ? 8'h8f : _GEN_882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_884 = 8'h74 == io_data_in[31:24] ? 8'h92 : _GEN_883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_885 = 8'h75 == io_data_in[31:24] ? 8'h9d : _GEN_884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_886 = 8'h76 == io_data_in[31:24] ? 8'h38 : _GEN_885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_887 = 8'h77 == io_data_in[31:24] ? 8'hf5 : _GEN_886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_888 = 8'h78 == io_data_in[31:24] ? 8'hbc : _GEN_887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_889 = 8'h79 == io_data_in[31:24] ? 8'hb6 : _GEN_888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_890 = 8'h7a == io_data_in[31:24] ? 8'hda : _GEN_889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_891 = 8'h7b == io_data_in[31:24] ? 8'h21 : _GEN_890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_892 = 8'h7c == io_data_in[31:24] ? 8'h10 : _GEN_891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_893 = 8'h7d == io_data_in[31:24] ? 8'hff : _GEN_892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_894 = 8'h7e == io_data_in[31:24] ? 8'hf3 : _GEN_893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_895 = 8'h7f == io_data_in[31:24] ? 8'hd2 : _GEN_894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_896 = 8'h80 == io_data_in[31:24] ? 8'hcd : _GEN_895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_897 = 8'h81 == io_data_in[31:24] ? 8'hc : _GEN_896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_898 = 8'h82 == io_data_in[31:24] ? 8'h13 : _GEN_897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_899 = 8'h83 == io_data_in[31:24] ? 8'hec : _GEN_898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_900 = 8'h84 == io_data_in[31:24] ? 8'h5f : _GEN_899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_901 = 8'h85 == io_data_in[31:24] ? 8'h97 : _GEN_900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_902 = 8'h86 == io_data_in[31:24] ? 8'h44 : _GEN_901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_903 = 8'h87 == io_data_in[31:24] ? 8'h17 : _GEN_902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_904 = 8'h88 == io_data_in[31:24] ? 8'hc4 : _GEN_903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_905 = 8'h89 == io_data_in[31:24] ? 8'ha7 : _GEN_904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_906 = 8'h8a == io_data_in[31:24] ? 8'h7e : _GEN_905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_907 = 8'h8b == io_data_in[31:24] ? 8'h3d : _GEN_906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_908 = 8'h8c == io_data_in[31:24] ? 8'h64 : _GEN_907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_909 = 8'h8d == io_data_in[31:24] ? 8'h5d : _GEN_908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_910 = 8'h8e == io_data_in[31:24] ? 8'h19 : _GEN_909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_911 = 8'h8f == io_data_in[31:24] ? 8'h73 : _GEN_910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_912 = 8'h90 == io_data_in[31:24] ? 8'h60 : _GEN_911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_913 = 8'h91 == io_data_in[31:24] ? 8'h81 : _GEN_912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_914 = 8'h92 == io_data_in[31:24] ? 8'h4f : _GEN_913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_915 = 8'h93 == io_data_in[31:24] ? 8'hdc : _GEN_914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_916 = 8'h94 == io_data_in[31:24] ? 8'h22 : _GEN_915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_917 = 8'h95 == io_data_in[31:24] ? 8'h2a : _GEN_916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_918 = 8'h96 == io_data_in[31:24] ? 8'h90 : _GEN_917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_919 = 8'h97 == io_data_in[31:24] ? 8'h88 : _GEN_918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_920 = 8'h98 == io_data_in[31:24] ? 8'h46 : _GEN_919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_921 = 8'h99 == io_data_in[31:24] ? 8'hee : _GEN_920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_922 = 8'h9a == io_data_in[31:24] ? 8'hb8 : _GEN_921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_923 = 8'h9b == io_data_in[31:24] ? 8'h14 : _GEN_922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_924 = 8'h9c == io_data_in[31:24] ? 8'hde : _GEN_923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_925 = 8'h9d == io_data_in[31:24] ? 8'h5e : _GEN_924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_926 = 8'h9e == io_data_in[31:24] ? 8'hb : _GEN_925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_927 = 8'h9f == io_data_in[31:24] ? 8'hdb : _GEN_926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_928 = 8'ha0 == io_data_in[31:24] ? 8'he0 : _GEN_927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_929 = 8'ha1 == io_data_in[31:24] ? 8'h32 : _GEN_928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_930 = 8'ha2 == io_data_in[31:24] ? 8'h3a : _GEN_929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_931 = 8'ha3 == io_data_in[31:24] ? 8'ha : _GEN_930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_932 = 8'ha4 == io_data_in[31:24] ? 8'h49 : _GEN_931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_933 = 8'ha5 == io_data_in[31:24] ? 8'h6 : _GEN_932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_934 = 8'ha6 == io_data_in[31:24] ? 8'h24 : _GEN_933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_935 = 8'ha7 == io_data_in[31:24] ? 8'h5c : _GEN_934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_936 = 8'ha8 == io_data_in[31:24] ? 8'hc2 : _GEN_935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_937 = 8'ha9 == io_data_in[31:24] ? 8'hd3 : _GEN_936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_938 = 8'haa == io_data_in[31:24] ? 8'hac : _GEN_937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_939 = 8'hab == io_data_in[31:24] ? 8'h62 : _GEN_938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_940 = 8'hac == io_data_in[31:24] ? 8'h91 : _GEN_939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_941 = 8'had == io_data_in[31:24] ? 8'h95 : _GEN_940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_942 = 8'hae == io_data_in[31:24] ? 8'he4 : _GEN_941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_943 = 8'haf == io_data_in[31:24] ? 8'h79 : _GEN_942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_944 = 8'hb0 == io_data_in[31:24] ? 8'he7 : _GEN_943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_945 = 8'hb1 == io_data_in[31:24] ? 8'hc8 : _GEN_944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_946 = 8'hb2 == io_data_in[31:24] ? 8'h37 : _GEN_945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_947 = 8'hb3 == io_data_in[31:24] ? 8'h6d : _GEN_946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_948 = 8'hb4 == io_data_in[31:24] ? 8'h8d : _GEN_947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_949 = 8'hb5 == io_data_in[31:24] ? 8'hd5 : _GEN_948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_950 = 8'hb6 == io_data_in[31:24] ? 8'h4e : _GEN_949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_951 = 8'hb7 == io_data_in[31:24] ? 8'ha9 : _GEN_950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_952 = 8'hb8 == io_data_in[31:24] ? 8'h6c : _GEN_951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_953 = 8'hb9 == io_data_in[31:24] ? 8'h56 : _GEN_952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_954 = 8'hba == io_data_in[31:24] ? 8'hf4 : _GEN_953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_955 = 8'hbb == io_data_in[31:24] ? 8'hea : _GEN_954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_956 = 8'hbc == io_data_in[31:24] ? 8'h65 : _GEN_955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_957 = 8'hbd == io_data_in[31:24] ? 8'h7a : _GEN_956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_958 = 8'hbe == io_data_in[31:24] ? 8'hae : _GEN_957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_959 = 8'hbf == io_data_in[31:24] ? 8'h8 : _GEN_958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_960 = 8'hc0 == io_data_in[31:24] ? 8'hba : _GEN_959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_961 = 8'hc1 == io_data_in[31:24] ? 8'h78 : _GEN_960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_962 = 8'hc2 == io_data_in[31:24] ? 8'h25 : _GEN_961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_963 = 8'hc3 == io_data_in[31:24] ? 8'h2e : _GEN_962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_964 = 8'hc4 == io_data_in[31:24] ? 8'h1c : _GEN_963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_965 = 8'hc5 == io_data_in[31:24] ? 8'ha6 : _GEN_964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_966 = 8'hc6 == io_data_in[31:24] ? 8'hb4 : _GEN_965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_967 = 8'hc7 == io_data_in[31:24] ? 8'hc6 : _GEN_966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_968 = 8'hc8 == io_data_in[31:24] ? 8'he8 : _GEN_967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_969 = 8'hc9 == io_data_in[31:24] ? 8'hdd : _GEN_968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_970 = 8'hca == io_data_in[31:24] ? 8'h74 : _GEN_969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_971 = 8'hcb == io_data_in[31:24] ? 8'h1f : _GEN_970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_972 = 8'hcc == io_data_in[31:24] ? 8'h4b : _GEN_971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_973 = 8'hcd == io_data_in[31:24] ? 8'hbd : _GEN_972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_974 = 8'hce == io_data_in[31:24] ? 8'h8b : _GEN_973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_975 = 8'hcf == io_data_in[31:24] ? 8'h8a : _GEN_974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_976 = 8'hd0 == io_data_in[31:24] ? 8'h70 : _GEN_975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_977 = 8'hd1 == io_data_in[31:24] ? 8'h3e : _GEN_976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_978 = 8'hd2 == io_data_in[31:24] ? 8'hb5 : _GEN_977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_979 = 8'hd3 == io_data_in[31:24] ? 8'h66 : _GEN_978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_980 = 8'hd4 == io_data_in[31:24] ? 8'h48 : _GEN_979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_981 = 8'hd5 == io_data_in[31:24] ? 8'h3 : _GEN_980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_982 = 8'hd6 == io_data_in[31:24] ? 8'hf6 : _GEN_981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_983 = 8'hd7 == io_data_in[31:24] ? 8'he : _GEN_982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_984 = 8'hd8 == io_data_in[31:24] ? 8'h61 : _GEN_983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_985 = 8'hd9 == io_data_in[31:24] ? 8'h35 : _GEN_984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_986 = 8'hda == io_data_in[31:24] ? 8'h57 : _GEN_985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_987 = 8'hdb == io_data_in[31:24] ? 8'hb9 : _GEN_986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_988 = 8'hdc == io_data_in[31:24] ? 8'h86 : _GEN_987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_989 = 8'hdd == io_data_in[31:24] ? 8'hc1 : _GEN_988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_990 = 8'hde == io_data_in[31:24] ? 8'h1d : _GEN_989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_991 = 8'hdf == io_data_in[31:24] ? 8'h9e : _GEN_990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_992 = 8'he0 == io_data_in[31:24] ? 8'he1 : _GEN_991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_993 = 8'he1 == io_data_in[31:24] ? 8'hf8 : _GEN_992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_994 = 8'he2 == io_data_in[31:24] ? 8'h98 : _GEN_993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_995 = 8'he3 == io_data_in[31:24] ? 8'h11 : _GEN_994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_996 = 8'he4 == io_data_in[31:24] ? 8'h69 : _GEN_995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_997 = 8'he5 == io_data_in[31:24] ? 8'hd9 : _GEN_996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_998 = 8'he6 == io_data_in[31:24] ? 8'h8e : _GEN_997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_999 = 8'he7 == io_data_in[31:24] ? 8'h94 : _GEN_998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1000 = 8'he8 == io_data_in[31:24] ? 8'h9b : _GEN_999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1001 = 8'he9 == io_data_in[31:24] ? 8'h1e : _GEN_1000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1002 = 8'hea == io_data_in[31:24] ? 8'h87 : _GEN_1001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1003 = 8'heb == io_data_in[31:24] ? 8'he9 : _GEN_1002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1004 = 8'hec == io_data_in[31:24] ? 8'hce : _GEN_1003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1005 = 8'hed == io_data_in[31:24] ? 8'h55 : _GEN_1004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1006 = 8'hee == io_data_in[31:24] ? 8'h28 : _GEN_1005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1007 = 8'hef == io_data_in[31:24] ? 8'hdf : _GEN_1006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1008 = 8'hf0 == io_data_in[31:24] ? 8'h8c : _GEN_1007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1009 = 8'hf1 == io_data_in[31:24] ? 8'ha1 : _GEN_1008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1010 = 8'hf2 == io_data_in[31:24] ? 8'h89 : _GEN_1009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1011 = 8'hf3 == io_data_in[31:24] ? 8'hd : _GEN_1010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1012 = 8'hf4 == io_data_in[31:24] ? 8'hbf : _GEN_1011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1013 = 8'hf5 == io_data_in[31:24] ? 8'he6 : _GEN_1012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1014 = 8'hf6 == io_data_in[31:24] ? 8'h42 : _GEN_1013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1015 = 8'hf7 == io_data_in[31:24] ? 8'h68 : _GEN_1014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1016 = 8'hf8 == io_data_in[31:24] ? 8'h41 : _GEN_1015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1017 = 8'hf9 == io_data_in[31:24] ? 8'h99 : _GEN_1016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1018 = 8'hfa == io_data_in[31:24] ? 8'h2d : _GEN_1017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1019 = 8'hfb == io_data_in[31:24] ? 8'hf : _GEN_1018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1020 = 8'hfc == io_data_in[31:24] ? 8'hb0 : _GEN_1019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1021 = 8'hfd == io_data_in[31:24] ? 8'h54 : _GEN_1020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1022 = 8'hfe == io_data_in[31:24] ? 8'hbb : _GEN_1021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1023 = 8'hff == io_data_in[31:24] ? 8'h16 : _GEN_1022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [15:0] io_data_out_hi = {_GEN_767,_GEN_1023}; // @[Cat.scala 30:58]
  XOR8 io_data_out_a ( // @[XOR32.scala 35:19]
    .io_data_in_1(io_data_out_a_io_data_in_1),
    .io_data_in_2(io_data_out_a_io_data_in_2),
    .io_data_out(io_data_out_a_io_data_out)
  );
  assign io_data_out = {io_data_out_hi,io_data_out_lo}; // @[Cat.scala 30:58]
  assign io_data_out_a_io_data_in_1 = 8'hff == io_data_in[15:8] ? 8'h16 : _GEN_254; // @[XOR32.scala 36:20 XOR32.scala 36:20]
  assign io_data_out_a_io_data_in_2 = io_rc_in; // @[XOR32.scala 37:20]
endmodule
module XOR32(
  input  [31:0] io_data_in_1,
  input  [31:0] io_data_in_2,
  output [31:0] io_data_out
);
  assign io_data_out = io_data_in_1 ^ io_data_in_2; // @[XOR32.scala 5:31]
endmodule
*/
module ShiftRows(
  input  [127:0] io_data_in,
  output [127:0] io_data_out
);
  wire [7:0] io_data_out_hi_hi_hi_hi = io_data_in[95:88]; // @[ShiftRows.scala 9:32]
  wire [7:0] io_data_out_hi_hi_hi_lo = io_data_in[55:48]; // @[ShiftRows.scala 9:50]
  wire [7:0] io_data_out_hi_hi_lo_hi = io_data_in[15:8]; // @[ShiftRows.scala 9:68]
  wire [7:0] io_data_out_hi_hi_lo_lo = io_data_in[103:96]; // @[ShiftRows.scala 9:85]
  wire [7:0] io_data_out_hi_lo_hi_hi = io_data_in[63:56]; // @[ShiftRows.scala 9:104]
  wire [7:0] io_data_out_hi_lo_hi_lo = io_data_in[23:16]; // @[ShiftRows.scala 9:122]
  wire [7:0] io_data_out_hi_lo_lo_hi = io_data_in[111:104]; // @[ShiftRows.scala 9:140]
  wire [7:0] io_data_out_hi_lo_lo_lo = io_data_in[71:64]; // @[ShiftRows.scala 9:160]
  wire [7:0] io_data_out_lo_hi_hi_hi = io_data_in[31:24]; // @[ShiftRows.scala 9:178]
  wire [7:0] io_data_out_lo_hi_hi_lo = io_data_in[119:112]; // @[ShiftRows.scala 9:197]
  wire [7:0] io_data_out_lo_hi_lo_hi = io_data_in[79:72]; // @[ShiftRows.scala 9:217]
  wire [7:0] io_data_out_lo_hi_lo_lo = io_data_in[39:32]; // @[ShiftRows.scala 9:235]
  wire [7:0] io_data_out_lo_lo_hi_hi = io_data_in[127:120]; // @[ShiftRows.scala 9:253]
  wire [7:0] io_data_out_lo_lo_hi_lo = io_data_in[87:80]; // @[ShiftRows.scala 9:273]
  wire [7:0] io_data_out_lo_lo_lo_hi = io_data_in[47:40]; // @[ShiftRows.scala 9:291]
  wire [7:0] io_data_out_lo_lo_lo_lo = io_data_in[7:0]; // @[ShiftRows.scala 9:309]
  wire [63:0] io_data_out_lo = {io_data_out_lo_hi_hi_hi,io_data_out_lo_hi_hi_lo,io_data_out_lo_hi_lo_hi,
    io_data_out_lo_hi_lo_lo,io_data_out_lo_lo_hi_hi,io_data_out_lo_lo_hi_lo,io_data_out_lo_lo_lo_hi,
    io_data_out_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] io_data_out_hi = {io_data_out_hi_hi_hi_hi,io_data_out_hi_hi_hi_lo,io_data_out_hi_hi_lo_hi,
    io_data_out_hi_hi_lo_lo,io_data_out_hi_lo_hi_hi,io_data_out_hi_lo_hi_lo,io_data_out_hi_lo_lo_hi,
    io_data_out_hi_lo_lo_lo}; // @[Cat.scala 30:58]
  assign io_data_out = {io_data_out_hi,io_data_out_lo}; // @[Cat.scala 30:58]
endmodule
module BS(
  input  [127:0] io_data_in,
  output [127:0] io_data_out
);
  wire [7:0] _GEN_1 = 8'h1 == io_data_in[15:8] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2 = 8'h2 == io_data_in[15:8] ? 8'h77 : _GEN_1; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3 = 8'h3 == io_data_in[15:8] ? 8'h7b : _GEN_2; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4 = 8'h4 == io_data_in[15:8] ? 8'hf2 : _GEN_3; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5 = 8'h5 == io_data_in[15:8] ? 8'h6b : _GEN_4; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6 = 8'h6 == io_data_in[15:8] ? 8'h6f : _GEN_5; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7 = 8'h7 == io_data_in[15:8] ? 8'hc5 : _GEN_6; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8 = 8'h8 == io_data_in[15:8] ? 8'h30 : _GEN_7; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9 = 8'h9 == io_data_in[15:8] ? 8'h1 : _GEN_8; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10 = 8'ha == io_data_in[15:8] ? 8'h67 : _GEN_9; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11 = 8'hb == io_data_in[15:8] ? 8'h2b : _GEN_10; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12 = 8'hc == io_data_in[15:8] ? 8'hfe : _GEN_11; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_13 = 8'hd == io_data_in[15:8] ? 8'hd7 : _GEN_12; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_14 = 8'he == io_data_in[15:8] ? 8'hab : _GEN_13; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_15 = 8'hf == io_data_in[15:8] ? 8'h76 : _GEN_14; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_16 = 8'h10 == io_data_in[15:8] ? 8'hca : _GEN_15; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_17 = 8'h11 == io_data_in[15:8] ? 8'h82 : _GEN_16; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_18 = 8'h12 == io_data_in[15:8] ? 8'hc9 : _GEN_17; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_19 = 8'h13 == io_data_in[15:8] ? 8'h7d : _GEN_18; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_20 = 8'h14 == io_data_in[15:8] ? 8'hfa : _GEN_19; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_21 = 8'h15 == io_data_in[15:8] ? 8'h59 : _GEN_20; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_22 = 8'h16 == io_data_in[15:8] ? 8'h47 : _GEN_21; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_23 = 8'h17 == io_data_in[15:8] ? 8'hf0 : _GEN_22; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_24 = 8'h18 == io_data_in[15:8] ? 8'had : _GEN_23; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_25 = 8'h19 == io_data_in[15:8] ? 8'hd4 : _GEN_24; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_26 = 8'h1a == io_data_in[15:8] ? 8'ha2 : _GEN_25; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_27 = 8'h1b == io_data_in[15:8] ? 8'haf : _GEN_26; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_28 = 8'h1c == io_data_in[15:8] ? 8'h9c : _GEN_27; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_29 = 8'h1d == io_data_in[15:8] ? 8'ha4 : _GEN_28; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_30 = 8'h1e == io_data_in[15:8] ? 8'h72 : _GEN_29; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_31 = 8'h1f == io_data_in[15:8] ? 8'hc0 : _GEN_30; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_32 = 8'h20 == io_data_in[15:8] ? 8'hb7 : _GEN_31; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_33 = 8'h21 == io_data_in[15:8] ? 8'hfd : _GEN_32; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_34 = 8'h22 == io_data_in[15:8] ? 8'h93 : _GEN_33; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_35 = 8'h23 == io_data_in[15:8] ? 8'h26 : _GEN_34; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_36 = 8'h24 == io_data_in[15:8] ? 8'h36 : _GEN_35; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_37 = 8'h25 == io_data_in[15:8] ? 8'h3f : _GEN_36; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_38 = 8'h26 == io_data_in[15:8] ? 8'hf7 : _GEN_37; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_39 = 8'h27 == io_data_in[15:8] ? 8'hcc : _GEN_38; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_40 = 8'h28 == io_data_in[15:8] ? 8'h34 : _GEN_39; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_41 = 8'h29 == io_data_in[15:8] ? 8'ha5 : _GEN_40; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_42 = 8'h2a == io_data_in[15:8] ? 8'he5 : _GEN_41; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_43 = 8'h2b == io_data_in[15:8] ? 8'hf1 : _GEN_42; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_44 = 8'h2c == io_data_in[15:8] ? 8'h71 : _GEN_43; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_45 = 8'h2d == io_data_in[15:8] ? 8'hd8 : _GEN_44; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_46 = 8'h2e == io_data_in[15:8] ? 8'h31 : _GEN_45; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_47 = 8'h2f == io_data_in[15:8] ? 8'h15 : _GEN_46; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_48 = 8'h30 == io_data_in[15:8] ? 8'h4 : _GEN_47; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_49 = 8'h31 == io_data_in[15:8] ? 8'hc7 : _GEN_48; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_50 = 8'h32 == io_data_in[15:8] ? 8'h23 : _GEN_49; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_51 = 8'h33 == io_data_in[15:8] ? 8'hc3 : _GEN_50; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_52 = 8'h34 == io_data_in[15:8] ? 8'h18 : _GEN_51; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_53 = 8'h35 == io_data_in[15:8] ? 8'h96 : _GEN_52; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_54 = 8'h36 == io_data_in[15:8] ? 8'h5 : _GEN_53; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_55 = 8'h37 == io_data_in[15:8] ? 8'h9a : _GEN_54; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_56 = 8'h38 == io_data_in[15:8] ? 8'h7 : _GEN_55; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_57 = 8'h39 == io_data_in[15:8] ? 8'h12 : _GEN_56; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_58 = 8'h3a == io_data_in[15:8] ? 8'h80 : _GEN_57; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_59 = 8'h3b == io_data_in[15:8] ? 8'he2 : _GEN_58; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_60 = 8'h3c == io_data_in[15:8] ? 8'heb : _GEN_59; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_61 = 8'h3d == io_data_in[15:8] ? 8'h27 : _GEN_60; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_62 = 8'h3e == io_data_in[15:8] ? 8'hb2 : _GEN_61; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_63 = 8'h3f == io_data_in[15:8] ? 8'h75 : _GEN_62; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_64 = 8'h40 == io_data_in[15:8] ? 8'h9 : _GEN_63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_65 = 8'h41 == io_data_in[15:8] ? 8'h83 : _GEN_64; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_66 = 8'h42 == io_data_in[15:8] ? 8'h2c : _GEN_65; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_67 = 8'h43 == io_data_in[15:8] ? 8'h1a : _GEN_66; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_68 = 8'h44 == io_data_in[15:8] ? 8'h1b : _GEN_67; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_69 = 8'h45 == io_data_in[15:8] ? 8'h6e : _GEN_68; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_70 = 8'h46 == io_data_in[15:8] ? 8'h5a : _GEN_69; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_71 = 8'h47 == io_data_in[15:8] ? 8'ha0 : _GEN_70; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_72 = 8'h48 == io_data_in[15:8] ? 8'h52 : _GEN_71; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_73 = 8'h49 == io_data_in[15:8] ? 8'h3b : _GEN_72; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_74 = 8'h4a == io_data_in[15:8] ? 8'hd6 : _GEN_73; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_75 = 8'h4b == io_data_in[15:8] ? 8'hb3 : _GEN_74; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_76 = 8'h4c == io_data_in[15:8] ? 8'h29 : _GEN_75; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_77 = 8'h4d == io_data_in[15:8] ? 8'he3 : _GEN_76; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_78 = 8'h4e == io_data_in[15:8] ? 8'h2f : _GEN_77; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_79 = 8'h4f == io_data_in[15:8] ? 8'h84 : _GEN_78; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_80 = 8'h50 == io_data_in[15:8] ? 8'h53 : _GEN_79; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_81 = 8'h51 == io_data_in[15:8] ? 8'hd1 : _GEN_80; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_82 = 8'h52 == io_data_in[15:8] ? 8'h0 : _GEN_81; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_83 = 8'h53 == io_data_in[15:8] ? 8'hed : _GEN_82; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_84 = 8'h54 == io_data_in[15:8] ? 8'h20 : _GEN_83; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_85 = 8'h55 == io_data_in[15:8] ? 8'hfc : _GEN_84; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_86 = 8'h56 == io_data_in[15:8] ? 8'hb1 : _GEN_85; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_87 = 8'h57 == io_data_in[15:8] ? 8'h5b : _GEN_86; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_88 = 8'h58 == io_data_in[15:8] ? 8'h6a : _GEN_87; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_89 = 8'h59 == io_data_in[15:8] ? 8'hcb : _GEN_88; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_90 = 8'h5a == io_data_in[15:8] ? 8'hbe : _GEN_89; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_91 = 8'h5b == io_data_in[15:8] ? 8'h39 : _GEN_90; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_92 = 8'h5c == io_data_in[15:8] ? 8'h4a : _GEN_91; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_93 = 8'h5d == io_data_in[15:8] ? 8'h4c : _GEN_92; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_94 = 8'h5e == io_data_in[15:8] ? 8'h58 : _GEN_93; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_95 = 8'h5f == io_data_in[15:8] ? 8'hcf : _GEN_94; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_96 = 8'h60 == io_data_in[15:8] ? 8'hd0 : _GEN_95; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_97 = 8'h61 == io_data_in[15:8] ? 8'hef : _GEN_96; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_98 = 8'h62 == io_data_in[15:8] ? 8'haa : _GEN_97; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_99 = 8'h63 == io_data_in[15:8] ? 8'hfb : _GEN_98; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_100 = 8'h64 == io_data_in[15:8] ? 8'h43 : _GEN_99; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_101 = 8'h65 == io_data_in[15:8] ? 8'h4d : _GEN_100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_102 = 8'h66 == io_data_in[15:8] ? 8'h33 : _GEN_101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_103 = 8'h67 == io_data_in[15:8] ? 8'h85 : _GEN_102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_104 = 8'h68 == io_data_in[15:8] ? 8'h45 : _GEN_103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_105 = 8'h69 == io_data_in[15:8] ? 8'hf9 : _GEN_104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_106 = 8'h6a == io_data_in[15:8] ? 8'h2 : _GEN_105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_107 = 8'h6b == io_data_in[15:8] ? 8'h7f : _GEN_106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_108 = 8'h6c == io_data_in[15:8] ? 8'h50 : _GEN_107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_109 = 8'h6d == io_data_in[15:8] ? 8'h3c : _GEN_108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_110 = 8'h6e == io_data_in[15:8] ? 8'h9f : _GEN_109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_111 = 8'h6f == io_data_in[15:8] ? 8'ha8 : _GEN_110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_112 = 8'h70 == io_data_in[15:8] ? 8'h51 : _GEN_111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_113 = 8'h71 == io_data_in[15:8] ? 8'ha3 : _GEN_112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_114 = 8'h72 == io_data_in[15:8] ? 8'h40 : _GEN_113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_115 = 8'h73 == io_data_in[15:8] ? 8'h8f : _GEN_114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_116 = 8'h74 == io_data_in[15:8] ? 8'h92 : _GEN_115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_117 = 8'h75 == io_data_in[15:8] ? 8'h9d : _GEN_116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_118 = 8'h76 == io_data_in[15:8] ? 8'h38 : _GEN_117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_119 = 8'h77 == io_data_in[15:8] ? 8'hf5 : _GEN_118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_120 = 8'h78 == io_data_in[15:8] ? 8'hbc : _GEN_119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_121 = 8'h79 == io_data_in[15:8] ? 8'hb6 : _GEN_120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_122 = 8'h7a == io_data_in[15:8] ? 8'hda : _GEN_121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_123 = 8'h7b == io_data_in[15:8] ? 8'h21 : _GEN_122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_124 = 8'h7c == io_data_in[15:8] ? 8'h10 : _GEN_123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_125 = 8'h7d == io_data_in[15:8] ? 8'hff : _GEN_124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_126 = 8'h7e == io_data_in[15:8] ? 8'hf3 : _GEN_125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_127 = 8'h7f == io_data_in[15:8] ? 8'hd2 : _GEN_126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_128 = 8'h80 == io_data_in[15:8] ? 8'hcd : _GEN_127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_129 = 8'h81 == io_data_in[15:8] ? 8'hc : _GEN_128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_130 = 8'h82 == io_data_in[15:8] ? 8'h13 : _GEN_129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_131 = 8'h83 == io_data_in[15:8] ? 8'hec : _GEN_130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_132 = 8'h84 == io_data_in[15:8] ? 8'h5f : _GEN_131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_133 = 8'h85 == io_data_in[15:8] ? 8'h97 : _GEN_132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_134 = 8'h86 == io_data_in[15:8] ? 8'h44 : _GEN_133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_135 = 8'h87 == io_data_in[15:8] ? 8'h17 : _GEN_134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_136 = 8'h88 == io_data_in[15:8] ? 8'hc4 : _GEN_135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_137 = 8'h89 == io_data_in[15:8] ? 8'ha7 : _GEN_136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_138 = 8'h8a == io_data_in[15:8] ? 8'h7e : _GEN_137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_139 = 8'h8b == io_data_in[15:8] ? 8'h3d : _GEN_138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_140 = 8'h8c == io_data_in[15:8] ? 8'h64 : _GEN_139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_141 = 8'h8d == io_data_in[15:8] ? 8'h5d : _GEN_140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_142 = 8'h8e == io_data_in[15:8] ? 8'h19 : _GEN_141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_143 = 8'h8f == io_data_in[15:8] ? 8'h73 : _GEN_142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_144 = 8'h90 == io_data_in[15:8] ? 8'h60 : _GEN_143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_145 = 8'h91 == io_data_in[15:8] ? 8'h81 : _GEN_144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_146 = 8'h92 == io_data_in[15:8] ? 8'h4f : _GEN_145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_147 = 8'h93 == io_data_in[15:8] ? 8'hdc : _GEN_146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_148 = 8'h94 == io_data_in[15:8] ? 8'h22 : _GEN_147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_149 = 8'h95 == io_data_in[15:8] ? 8'h2a : _GEN_148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_150 = 8'h96 == io_data_in[15:8] ? 8'h90 : _GEN_149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_151 = 8'h97 == io_data_in[15:8] ? 8'h88 : _GEN_150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_152 = 8'h98 == io_data_in[15:8] ? 8'h46 : _GEN_151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_153 = 8'h99 == io_data_in[15:8] ? 8'hee : _GEN_152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_154 = 8'h9a == io_data_in[15:8] ? 8'hb8 : _GEN_153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_155 = 8'h9b == io_data_in[15:8] ? 8'h14 : _GEN_154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_156 = 8'h9c == io_data_in[15:8] ? 8'hde : _GEN_155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_157 = 8'h9d == io_data_in[15:8] ? 8'h5e : _GEN_156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_158 = 8'h9e == io_data_in[15:8] ? 8'hb : _GEN_157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_159 = 8'h9f == io_data_in[15:8] ? 8'hdb : _GEN_158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_160 = 8'ha0 == io_data_in[15:8] ? 8'he0 : _GEN_159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_161 = 8'ha1 == io_data_in[15:8] ? 8'h32 : _GEN_160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_162 = 8'ha2 == io_data_in[15:8] ? 8'h3a : _GEN_161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_163 = 8'ha3 == io_data_in[15:8] ? 8'ha : _GEN_162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_164 = 8'ha4 == io_data_in[15:8] ? 8'h49 : _GEN_163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_165 = 8'ha5 == io_data_in[15:8] ? 8'h6 : _GEN_164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_166 = 8'ha6 == io_data_in[15:8] ? 8'h24 : _GEN_165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_167 = 8'ha7 == io_data_in[15:8] ? 8'h5c : _GEN_166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_168 = 8'ha8 == io_data_in[15:8] ? 8'hc2 : _GEN_167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_169 = 8'ha9 == io_data_in[15:8] ? 8'hd3 : _GEN_168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_170 = 8'haa == io_data_in[15:8] ? 8'hac : _GEN_169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_171 = 8'hab == io_data_in[15:8] ? 8'h62 : _GEN_170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_172 = 8'hac == io_data_in[15:8] ? 8'h91 : _GEN_171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_173 = 8'had == io_data_in[15:8] ? 8'h95 : _GEN_172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_174 = 8'hae == io_data_in[15:8] ? 8'he4 : _GEN_173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_175 = 8'haf == io_data_in[15:8] ? 8'h79 : _GEN_174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_176 = 8'hb0 == io_data_in[15:8] ? 8'he7 : _GEN_175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_177 = 8'hb1 == io_data_in[15:8] ? 8'hc8 : _GEN_176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_178 = 8'hb2 == io_data_in[15:8] ? 8'h37 : _GEN_177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_179 = 8'hb3 == io_data_in[15:8] ? 8'h6d : _GEN_178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_180 = 8'hb4 == io_data_in[15:8] ? 8'h8d : _GEN_179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_181 = 8'hb5 == io_data_in[15:8] ? 8'hd5 : _GEN_180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_182 = 8'hb6 == io_data_in[15:8] ? 8'h4e : _GEN_181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_183 = 8'hb7 == io_data_in[15:8] ? 8'ha9 : _GEN_182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_184 = 8'hb8 == io_data_in[15:8] ? 8'h6c : _GEN_183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_185 = 8'hb9 == io_data_in[15:8] ? 8'h56 : _GEN_184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_186 = 8'hba == io_data_in[15:8] ? 8'hf4 : _GEN_185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_187 = 8'hbb == io_data_in[15:8] ? 8'hea : _GEN_186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_188 = 8'hbc == io_data_in[15:8] ? 8'h65 : _GEN_187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_189 = 8'hbd == io_data_in[15:8] ? 8'h7a : _GEN_188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_190 = 8'hbe == io_data_in[15:8] ? 8'hae : _GEN_189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_191 = 8'hbf == io_data_in[15:8] ? 8'h8 : _GEN_190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_192 = 8'hc0 == io_data_in[15:8] ? 8'hba : _GEN_191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_193 = 8'hc1 == io_data_in[15:8] ? 8'h78 : _GEN_192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_194 = 8'hc2 == io_data_in[15:8] ? 8'h25 : _GEN_193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_195 = 8'hc3 == io_data_in[15:8] ? 8'h2e : _GEN_194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_196 = 8'hc4 == io_data_in[15:8] ? 8'h1c : _GEN_195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_197 = 8'hc5 == io_data_in[15:8] ? 8'ha6 : _GEN_196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_198 = 8'hc6 == io_data_in[15:8] ? 8'hb4 : _GEN_197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_199 = 8'hc7 == io_data_in[15:8] ? 8'hc6 : _GEN_198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_200 = 8'hc8 == io_data_in[15:8] ? 8'he8 : _GEN_199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_201 = 8'hc9 == io_data_in[15:8] ? 8'hdd : _GEN_200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_202 = 8'hca == io_data_in[15:8] ? 8'h74 : _GEN_201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_203 = 8'hcb == io_data_in[15:8] ? 8'h1f : _GEN_202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_204 = 8'hcc == io_data_in[15:8] ? 8'h4b : _GEN_203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_205 = 8'hcd == io_data_in[15:8] ? 8'hbd : _GEN_204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_206 = 8'hce == io_data_in[15:8] ? 8'h8b : _GEN_205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_207 = 8'hcf == io_data_in[15:8] ? 8'h8a : _GEN_206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_208 = 8'hd0 == io_data_in[15:8] ? 8'h70 : _GEN_207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_209 = 8'hd1 == io_data_in[15:8] ? 8'h3e : _GEN_208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_210 = 8'hd2 == io_data_in[15:8] ? 8'hb5 : _GEN_209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_211 = 8'hd3 == io_data_in[15:8] ? 8'h66 : _GEN_210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_212 = 8'hd4 == io_data_in[15:8] ? 8'h48 : _GEN_211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_213 = 8'hd5 == io_data_in[15:8] ? 8'h3 : _GEN_212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_214 = 8'hd6 == io_data_in[15:8] ? 8'hf6 : _GEN_213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_215 = 8'hd7 == io_data_in[15:8] ? 8'he : _GEN_214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_216 = 8'hd8 == io_data_in[15:8] ? 8'h61 : _GEN_215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_217 = 8'hd9 == io_data_in[15:8] ? 8'h35 : _GEN_216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_218 = 8'hda == io_data_in[15:8] ? 8'h57 : _GEN_217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_219 = 8'hdb == io_data_in[15:8] ? 8'hb9 : _GEN_218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_220 = 8'hdc == io_data_in[15:8] ? 8'h86 : _GEN_219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_221 = 8'hdd == io_data_in[15:8] ? 8'hc1 : _GEN_220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_222 = 8'hde == io_data_in[15:8] ? 8'h1d : _GEN_221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_223 = 8'hdf == io_data_in[15:8] ? 8'h9e : _GEN_222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_224 = 8'he0 == io_data_in[15:8] ? 8'he1 : _GEN_223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_225 = 8'he1 == io_data_in[15:8] ? 8'hf8 : _GEN_224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_226 = 8'he2 == io_data_in[15:8] ? 8'h98 : _GEN_225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_227 = 8'he3 == io_data_in[15:8] ? 8'h11 : _GEN_226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_228 = 8'he4 == io_data_in[15:8] ? 8'h69 : _GEN_227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_229 = 8'he5 == io_data_in[15:8] ? 8'hd9 : _GEN_228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_230 = 8'he6 == io_data_in[15:8] ? 8'h8e : _GEN_229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_231 = 8'he7 == io_data_in[15:8] ? 8'h94 : _GEN_230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_232 = 8'he8 == io_data_in[15:8] ? 8'h9b : _GEN_231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_233 = 8'he9 == io_data_in[15:8] ? 8'h1e : _GEN_232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_234 = 8'hea == io_data_in[15:8] ? 8'h87 : _GEN_233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_235 = 8'heb == io_data_in[15:8] ? 8'he9 : _GEN_234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_236 = 8'hec == io_data_in[15:8] ? 8'hce : _GEN_235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_237 = 8'hed == io_data_in[15:8] ? 8'h55 : _GEN_236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_238 = 8'hee == io_data_in[15:8] ? 8'h28 : _GEN_237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_239 = 8'hef == io_data_in[15:8] ? 8'hdf : _GEN_238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_240 = 8'hf0 == io_data_in[15:8] ? 8'h8c : _GEN_239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_241 = 8'hf1 == io_data_in[15:8] ? 8'ha1 : _GEN_240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_242 = 8'hf2 == io_data_in[15:8] ? 8'h89 : _GEN_241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_243 = 8'hf3 == io_data_in[15:8] ? 8'hd : _GEN_242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_244 = 8'hf4 == io_data_in[15:8] ? 8'hbf : _GEN_243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_245 = 8'hf5 == io_data_in[15:8] ? 8'he6 : _GEN_244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_246 = 8'hf6 == io_data_in[15:8] ? 8'h42 : _GEN_245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_247 = 8'hf7 == io_data_in[15:8] ? 8'h68 : _GEN_246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_248 = 8'hf8 == io_data_in[15:8] ? 8'h41 : _GEN_247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_249 = 8'hf9 == io_data_in[15:8] ? 8'h99 : _GEN_248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_250 = 8'hfa == io_data_in[15:8] ? 8'h2d : _GEN_249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_251 = 8'hfb == io_data_in[15:8] ? 8'hf : _GEN_250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_252 = 8'hfc == io_data_in[15:8] ? 8'hb0 : _GEN_251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_253 = 8'hfd == io_data_in[15:8] ? 8'h54 : _GEN_252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_254 = 8'hfe == io_data_in[15:8] ? 8'hbb : _GEN_253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_255 = 8'hff == io_data_in[15:8] ? 8'h16 : _GEN_254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_257 = 8'h1 == io_data_in[7:0] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_258 = 8'h2 == io_data_in[7:0] ? 8'h77 : _GEN_257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_259 = 8'h3 == io_data_in[7:0] ? 8'h7b : _GEN_258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_260 = 8'h4 == io_data_in[7:0] ? 8'hf2 : _GEN_259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_261 = 8'h5 == io_data_in[7:0] ? 8'h6b : _GEN_260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_262 = 8'h6 == io_data_in[7:0] ? 8'h6f : _GEN_261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_263 = 8'h7 == io_data_in[7:0] ? 8'hc5 : _GEN_262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_264 = 8'h8 == io_data_in[7:0] ? 8'h30 : _GEN_263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_265 = 8'h9 == io_data_in[7:0] ? 8'h1 : _GEN_264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_266 = 8'ha == io_data_in[7:0] ? 8'h67 : _GEN_265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_267 = 8'hb == io_data_in[7:0] ? 8'h2b : _GEN_266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_268 = 8'hc == io_data_in[7:0] ? 8'hfe : _GEN_267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_269 = 8'hd == io_data_in[7:0] ? 8'hd7 : _GEN_268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_270 = 8'he == io_data_in[7:0] ? 8'hab : _GEN_269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_271 = 8'hf == io_data_in[7:0] ? 8'h76 : _GEN_270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_272 = 8'h10 == io_data_in[7:0] ? 8'hca : _GEN_271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_273 = 8'h11 == io_data_in[7:0] ? 8'h82 : _GEN_272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_274 = 8'h12 == io_data_in[7:0] ? 8'hc9 : _GEN_273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_275 = 8'h13 == io_data_in[7:0] ? 8'h7d : _GEN_274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_276 = 8'h14 == io_data_in[7:0] ? 8'hfa : _GEN_275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_277 = 8'h15 == io_data_in[7:0] ? 8'h59 : _GEN_276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_278 = 8'h16 == io_data_in[7:0] ? 8'h47 : _GEN_277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_279 = 8'h17 == io_data_in[7:0] ? 8'hf0 : _GEN_278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_280 = 8'h18 == io_data_in[7:0] ? 8'had : _GEN_279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_281 = 8'h19 == io_data_in[7:0] ? 8'hd4 : _GEN_280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_282 = 8'h1a == io_data_in[7:0] ? 8'ha2 : _GEN_281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_283 = 8'h1b == io_data_in[7:0] ? 8'haf : _GEN_282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_284 = 8'h1c == io_data_in[7:0] ? 8'h9c : _GEN_283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_285 = 8'h1d == io_data_in[7:0] ? 8'ha4 : _GEN_284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_286 = 8'h1e == io_data_in[7:0] ? 8'h72 : _GEN_285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_287 = 8'h1f == io_data_in[7:0] ? 8'hc0 : _GEN_286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_288 = 8'h20 == io_data_in[7:0] ? 8'hb7 : _GEN_287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_289 = 8'h21 == io_data_in[7:0] ? 8'hfd : _GEN_288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_290 = 8'h22 == io_data_in[7:0] ? 8'h93 : _GEN_289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_291 = 8'h23 == io_data_in[7:0] ? 8'h26 : _GEN_290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_292 = 8'h24 == io_data_in[7:0] ? 8'h36 : _GEN_291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_293 = 8'h25 == io_data_in[7:0] ? 8'h3f : _GEN_292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_294 = 8'h26 == io_data_in[7:0] ? 8'hf7 : _GEN_293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_295 = 8'h27 == io_data_in[7:0] ? 8'hcc : _GEN_294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_296 = 8'h28 == io_data_in[7:0] ? 8'h34 : _GEN_295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_297 = 8'h29 == io_data_in[7:0] ? 8'ha5 : _GEN_296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_298 = 8'h2a == io_data_in[7:0] ? 8'he5 : _GEN_297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_299 = 8'h2b == io_data_in[7:0] ? 8'hf1 : _GEN_298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_300 = 8'h2c == io_data_in[7:0] ? 8'h71 : _GEN_299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_301 = 8'h2d == io_data_in[7:0] ? 8'hd8 : _GEN_300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_302 = 8'h2e == io_data_in[7:0] ? 8'h31 : _GEN_301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_303 = 8'h2f == io_data_in[7:0] ? 8'h15 : _GEN_302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_304 = 8'h30 == io_data_in[7:0] ? 8'h4 : _GEN_303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_305 = 8'h31 == io_data_in[7:0] ? 8'hc7 : _GEN_304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_306 = 8'h32 == io_data_in[7:0] ? 8'h23 : _GEN_305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_307 = 8'h33 == io_data_in[7:0] ? 8'hc3 : _GEN_306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_308 = 8'h34 == io_data_in[7:0] ? 8'h18 : _GEN_307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_309 = 8'h35 == io_data_in[7:0] ? 8'h96 : _GEN_308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_310 = 8'h36 == io_data_in[7:0] ? 8'h5 : _GEN_309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_311 = 8'h37 == io_data_in[7:0] ? 8'h9a : _GEN_310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_312 = 8'h38 == io_data_in[7:0] ? 8'h7 : _GEN_311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_313 = 8'h39 == io_data_in[7:0] ? 8'h12 : _GEN_312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_314 = 8'h3a == io_data_in[7:0] ? 8'h80 : _GEN_313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_315 = 8'h3b == io_data_in[7:0] ? 8'he2 : _GEN_314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_316 = 8'h3c == io_data_in[7:0] ? 8'heb : _GEN_315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_317 = 8'h3d == io_data_in[7:0] ? 8'h27 : _GEN_316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_318 = 8'h3e == io_data_in[7:0] ? 8'hb2 : _GEN_317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_319 = 8'h3f == io_data_in[7:0] ? 8'h75 : _GEN_318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_320 = 8'h40 == io_data_in[7:0] ? 8'h9 : _GEN_319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_321 = 8'h41 == io_data_in[7:0] ? 8'h83 : _GEN_320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_322 = 8'h42 == io_data_in[7:0] ? 8'h2c : _GEN_321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_323 = 8'h43 == io_data_in[7:0] ? 8'h1a : _GEN_322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_324 = 8'h44 == io_data_in[7:0] ? 8'h1b : _GEN_323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_325 = 8'h45 == io_data_in[7:0] ? 8'h6e : _GEN_324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_326 = 8'h46 == io_data_in[7:0] ? 8'h5a : _GEN_325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_327 = 8'h47 == io_data_in[7:0] ? 8'ha0 : _GEN_326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_328 = 8'h48 == io_data_in[7:0] ? 8'h52 : _GEN_327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_329 = 8'h49 == io_data_in[7:0] ? 8'h3b : _GEN_328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_330 = 8'h4a == io_data_in[7:0] ? 8'hd6 : _GEN_329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_331 = 8'h4b == io_data_in[7:0] ? 8'hb3 : _GEN_330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_332 = 8'h4c == io_data_in[7:0] ? 8'h29 : _GEN_331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_333 = 8'h4d == io_data_in[7:0] ? 8'he3 : _GEN_332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_334 = 8'h4e == io_data_in[7:0] ? 8'h2f : _GEN_333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_335 = 8'h4f == io_data_in[7:0] ? 8'h84 : _GEN_334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_336 = 8'h50 == io_data_in[7:0] ? 8'h53 : _GEN_335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_337 = 8'h51 == io_data_in[7:0] ? 8'hd1 : _GEN_336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_338 = 8'h52 == io_data_in[7:0] ? 8'h0 : _GEN_337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_339 = 8'h53 == io_data_in[7:0] ? 8'hed : _GEN_338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_340 = 8'h54 == io_data_in[7:0] ? 8'h20 : _GEN_339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_341 = 8'h55 == io_data_in[7:0] ? 8'hfc : _GEN_340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_342 = 8'h56 == io_data_in[7:0] ? 8'hb1 : _GEN_341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_343 = 8'h57 == io_data_in[7:0] ? 8'h5b : _GEN_342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_344 = 8'h58 == io_data_in[7:0] ? 8'h6a : _GEN_343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_345 = 8'h59 == io_data_in[7:0] ? 8'hcb : _GEN_344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_346 = 8'h5a == io_data_in[7:0] ? 8'hbe : _GEN_345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_347 = 8'h5b == io_data_in[7:0] ? 8'h39 : _GEN_346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_348 = 8'h5c == io_data_in[7:0] ? 8'h4a : _GEN_347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_349 = 8'h5d == io_data_in[7:0] ? 8'h4c : _GEN_348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_350 = 8'h5e == io_data_in[7:0] ? 8'h58 : _GEN_349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_351 = 8'h5f == io_data_in[7:0] ? 8'hcf : _GEN_350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_352 = 8'h60 == io_data_in[7:0] ? 8'hd0 : _GEN_351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_353 = 8'h61 == io_data_in[7:0] ? 8'hef : _GEN_352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_354 = 8'h62 == io_data_in[7:0] ? 8'haa : _GEN_353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_355 = 8'h63 == io_data_in[7:0] ? 8'hfb : _GEN_354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_356 = 8'h64 == io_data_in[7:0] ? 8'h43 : _GEN_355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_357 = 8'h65 == io_data_in[7:0] ? 8'h4d : _GEN_356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_358 = 8'h66 == io_data_in[7:0] ? 8'h33 : _GEN_357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_359 = 8'h67 == io_data_in[7:0] ? 8'h85 : _GEN_358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_360 = 8'h68 == io_data_in[7:0] ? 8'h45 : _GEN_359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_361 = 8'h69 == io_data_in[7:0] ? 8'hf9 : _GEN_360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_362 = 8'h6a == io_data_in[7:0] ? 8'h2 : _GEN_361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_363 = 8'h6b == io_data_in[7:0] ? 8'h7f : _GEN_362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_364 = 8'h6c == io_data_in[7:0] ? 8'h50 : _GEN_363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_365 = 8'h6d == io_data_in[7:0] ? 8'h3c : _GEN_364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_366 = 8'h6e == io_data_in[7:0] ? 8'h9f : _GEN_365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_367 = 8'h6f == io_data_in[7:0] ? 8'ha8 : _GEN_366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_368 = 8'h70 == io_data_in[7:0] ? 8'h51 : _GEN_367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_369 = 8'h71 == io_data_in[7:0] ? 8'ha3 : _GEN_368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_370 = 8'h72 == io_data_in[7:0] ? 8'h40 : _GEN_369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_371 = 8'h73 == io_data_in[7:0] ? 8'h8f : _GEN_370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_372 = 8'h74 == io_data_in[7:0] ? 8'h92 : _GEN_371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_373 = 8'h75 == io_data_in[7:0] ? 8'h9d : _GEN_372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_374 = 8'h76 == io_data_in[7:0] ? 8'h38 : _GEN_373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_375 = 8'h77 == io_data_in[7:0] ? 8'hf5 : _GEN_374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_376 = 8'h78 == io_data_in[7:0] ? 8'hbc : _GEN_375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_377 = 8'h79 == io_data_in[7:0] ? 8'hb6 : _GEN_376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_378 = 8'h7a == io_data_in[7:0] ? 8'hda : _GEN_377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_379 = 8'h7b == io_data_in[7:0] ? 8'h21 : _GEN_378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_380 = 8'h7c == io_data_in[7:0] ? 8'h10 : _GEN_379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_381 = 8'h7d == io_data_in[7:0] ? 8'hff : _GEN_380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_382 = 8'h7e == io_data_in[7:0] ? 8'hf3 : _GEN_381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_383 = 8'h7f == io_data_in[7:0] ? 8'hd2 : _GEN_382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_384 = 8'h80 == io_data_in[7:0] ? 8'hcd : _GEN_383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_385 = 8'h81 == io_data_in[7:0] ? 8'hc : _GEN_384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_386 = 8'h82 == io_data_in[7:0] ? 8'h13 : _GEN_385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_387 = 8'h83 == io_data_in[7:0] ? 8'hec : _GEN_386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_388 = 8'h84 == io_data_in[7:0] ? 8'h5f : _GEN_387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_389 = 8'h85 == io_data_in[7:0] ? 8'h97 : _GEN_388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_390 = 8'h86 == io_data_in[7:0] ? 8'h44 : _GEN_389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_391 = 8'h87 == io_data_in[7:0] ? 8'h17 : _GEN_390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_392 = 8'h88 == io_data_in[7:0] ? 8'hc4 : _GEN_391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_393 = 8'h89 == io_data_in[7:0] ? 8'ha7 : _GEN_392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_394 = 8'h8a == io_data_in[7:0] ? 8'h7e : _GEN_393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_395 = 8'h8b == io_data_in[7:0] ? 8'h3d : _GEN_394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_396 = 8'h8c == io_data_in[7:0] ? 8'h64 : _GEN_395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_397 = 8'h8d == io_data_in[7:0] ? 8'h5d : _GEN_396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_398 = 8'h8e == io_data_in[7:0] ? 8'h19 : _GEN_397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_399 = 8'h8f == io_data_in[7:0] ? 8'h73 : _GEN_398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_400 = 8'h90 == io_data_in[7:0] ? 8'h60 : _GEN_399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_401 = 8'h91 == io_data_in[7:0] ? 8'h81 : _GEN_400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_402 = 8'h92 == io_data_in[7:0] ? 8'h4f : _GEN_401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_403 = 8'h93 == io_data_in[7:0] ? 8'hdc : _GEN_402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_404 = 8'h94 == io_data_in[7:0] ? 8'h22 : _GEN_403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_405 = 8'h95 == io_data_in[7:0] ? 8'h2a : _GEN_404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_406 = 8'h96 == io_data_in[7:0] ? 8'h90 : _GEN_405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_407 = 8'h97 == io_data_in[7:0] ? 8'h88 : _GEN_406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_408 = 8'h98 == io_data_in[7:0] ? 8'h46 : _GEN_407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_409 = 8'h99 == io_data_in[7:0] ? 8'hee : _GEN_408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_410 = 8'h9a == io_data_in[7:0] ? 8'hb8 : _GEN_409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_411 = 8'h9b == io_data_in[7:0] ? 8'h14 : _GEN_410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_412 = 8'h9c == io_data_in[7:0] ? 8'hde : _GEN_411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_413 = 8'h9d == io_data_in[7:0] ? 8'h5e : _GEN_412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_414 = 8'h9e == io_data_in[7:0] ? 8'hb : _GEN_413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_415 = 8'h9f == io_data_in[7:0] ? 8'hdb : _GEN_414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_416 = 8'ha0 == io_data_in[7:0] ? 8'he0 : _GEN_415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_417 = 8'ha1 == io_data_in[7:0] ? 8'h32 : _GEN_416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_418 = 8'ha2 == io_data_in[7:0] ? 8'h3a : _GEN_417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_419 = 8'ha3 == io_data_in[7:0] ? 8'ha : _GEN_418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_420 = 8'ha4 == io_data_in[7:0] ? 8'h49 : _GEN_419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_421 = 8'ha5 == io_data_in[7:0] ? 8'h6 : _GEN_420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_422 = 8'ha6 == io_data_in[7:0] ? 8'h24 : _GEN_421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_423 = 8'ha7 == io_data_in[7:0] ? 8'h5c : _GEN_422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_424 = 8'ha8 == io_data_in[7:0] ? 8'hc2 : _GEN_423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_425 = 8'ha9 == io_data_in[7:0] ? 8'hd3 : _GEN_424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_426 = 8'haa == io_data_in[7:0] ? 8'hac : _GEN_425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_427 = 8'hab == io_data_in[7:0] ? 8'h62 : _GEN_426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_428 = 8'hac == io_data_in[7:0] ? 8'h91 : _GEN_427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_429 = 8'had == io_data_in[7:0] ? 8'h95 : _GEN_428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_430 = 8'hae == io_data_in[7:0] ? 8'he4 : _GEN_429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_431 = 8'haf == io_data_in[7:0] ? 8'h79 : _GEN_430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_432 = 8'hb0 == io_data_in[7:0] ? 8'he7 : _GEN_431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_433 = 8'hb1 == io_data_in[7:0] ? 8'hc8 : _GEN_432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_434 = 8'hb2 == io_data_in[7:0] ? 8'h37 : _GEN_433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_435 = 8'hb3 == io_data_in[7:0] ? 8'h6d : _GEN_434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_436 = 8'hb4 == io_data_in[7:0] ? 8'h8d : _GEN_435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_437 = 8'hb5 == io_data_in[7:0] ? 8'hd5 : _GEN_436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_438 = 8'hb6 == io_data_in[7:0] ? 8'h4e : _GEN_437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_439 = 8'hb7 == io_data_in[7:0] ? 8'ha9 : _GEN_438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_440 = 8'hb8 == io_data_in[7:0] ? 8'h6c : _GEN_439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_441 = 8'hb9 == io_data_in[7:0] ? 8'h56 : _GEN_440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_442 = 8'hba == io_data_in[7:0] ? 8'hf4 : _GEN_441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_443 = 8'hbb == io_data_in[7:0] ? 8'hea : _GEN_442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_444 = 8'hbc == io_data_in[7:0] ? 8'h65 : _GEN_443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_445 = 8'hbd == io_data_in[7:0] ? 8'h7a : _GEN_444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_446 = 8'hbe == io_data_in[7:0] ? 8'hae : _GEN_445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_447 = 8'hbf == io_data_in[7:0] ? 8'h8 : _GEN_446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_448 = 8'hc0 == io_data_in[7:0] ? 8'hba : _GEN_447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_449 = 8'hc1 == io_data_in[7:0] ? 8'h78 : _GEN_448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_450 = 8'hc2 == io_data_in[7:0] ? 8'h25 : _GEN_449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_451 = 8'hc3 == io_data_in[7:0] ? 8'h2e : _GEN_450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_452 = 8'hc4 == io_data_in[7:0] ? 8'h1c : _GEN_451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_453 = 8'hc5 == io_data_in[7:0] ? 8'ha6 : _GEN_452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_454 = 8'hc6 == io_data_in[7:0] ? 8'hb4 : _GEN_453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_455 = 8'hc7 == io_data_in[7:0] ? 8'hc6 : _GEN_454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_456 = 8'hc8 == io_data_in[7:0] ? 8'he8 : _GEN_455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_457 = 8'hc9 == io_data_in[7:0] ? 8'hdd : _GEN_456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_458 = 8'hca == io_data_in[7:0] ? 8'h74 : _GEN_457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_459 = 8'hcb == io_data_in[7:0] ? 8'h1f : _GEN_458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_460 = 8'hcc == io_data_in[7:0] ? 8'h4b : _GEN_459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_461 = 8'hcd == io_data_in[7:0] ? 8'hbd : _GEN_460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_462 = 8'hce == io_data_in[7:0] ? 8'h8b : _GEN_461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_463 = 8'hcf == io_data_in[7:0] ? 8'h8a : _GEN_462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_464 = 8'hd0 == io_data_in[7:0] ? 8'h70 : _GEN_463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_465 = 8'hd1 == io_data_in[7:0] ? 8'h3e : _GEN_464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_466 = 8'hd2 == io_data_in[7:0] ? 8'hb5 : _GEN_465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_467 = 8'hd3 == io_data_in[7:0] ? 8'h66 : _GEN_466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_468 = 8'hd4 == io_data_in[7:0] ? 8'h48 : _GEN_467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_469 = 8'hd5 == io_data_in[7:0] ? 8'h3 : _GEN_468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_470 = 8'hd6 == io_data_in[7:0] ? 8'hf6 : _GEN_469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_471 = 8'hd7 == io_data_in[7:0] ? 8'he : _GEN_470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_472 = 8'hd8 == io_data_in[7:0] ? 8'h61 : _GEN_471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_473 = 8'hd9 == io_data_in[7:0] ? 8'h35 : _GEN_472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_474 = 8'hda == io_data_in[7:0] ? 8'h57 : _GEN_473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_475 = 8'hdb == io_data_in[7:0] ? 8'hb9 : _GEN_474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_476 = 8'hdc == io_data_in[7:0] ? 8'h86 : _GEN_475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_477 = 8'hdd == io_data_in[7:0] ? 8'hc1 : _GEN_476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_478 = 8'hde == io_data_in[7:0] ? 8'h1d : _GEN_477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_479 = 8'hdf == io_data_in[7:0] ? 8'h9e : _GEN_478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_480 = 8'he0 == io_data_in[7:0] ? 8'he1 : _GEN_479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_481 = 8'he1 == io_data_in[7:0] ? 8'hf8 : _GEN_480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_482 = 8'he2 == io_data_in[7:0] ? 8'h98 : _GEN_481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_483 = 8'he3 == io_data_in[7:0] ? 8'h11 : _GEN_482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_484 = 8'he4 == io_data_in[7:0] ? 8'h69 : _GEN_483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_485 = 8'he5 == io_data_in[7:0] ? 8'hd9 : _GEN_484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_486 = 8'he6 == io_data_in[7:0] ? 8'h8e : _GEN_485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_487 = 8'he7 == io_data_in[7:0] ? 8'h94 : _GEN_486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_488 = 8'he8 == io_data_in[7:0] ? 8'h9b : _GEN_487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_489 = 8'he9 == io_data_in[7:0] ? 8'h1e : _GEN_488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_490 = 8'hea == io_data_in[7:0] ? 8'h87 : _GEN_489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_491 = 8'heb == io_data_in[7:0] ? 8'he9 : _GEN_490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_492 = 8'hec == io_data_in[7:0] ? 8'hce : _GEN_491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_493 = 8'hed == io_data_in[7:0] ? 8'h55 : _GEN_492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_494 = 8'hee == io_data_in[7:0] ? 8'h28 : _GEN_493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_495 = 8'hef == io_data_in[7:0] ? 8'hdf : _GEN_494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_496 = 8'hf0 == io_data_in[7:0] ? 8'h8c : _GEN_495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_497 = 8'hf1 == io_data_in[7:0] ? 8'ha1 : _GEN_496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_498 = 8'hf2 == io_data_in[7:0] ? 8'h89 : _GEN_497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_499 = 8'hf3 == io_data_in[7:0] ? 8'hd : _GEN_498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_500 = 8'hf4 == io_data_in[7:0] ? 8'hbf : _GEN_499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_501 = 8'hf5 == io_data_in[7:0] ? 8'he6 : _GEN_500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_502 = 8'hf6 == io_data_in[7:0] ? 8'h42 : _GEN_501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_503 = 8'hf7 == io_data_in[7:0] ? 8'h68 : _GEN_502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_504 = 8'hf8 == io_data_in[7:0] ? 8'h41 : _GEN_503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_505 = 8'hf9 == io_data_in[7:0] ? 8'h99 : _GEN_504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_506 = 8'hfa == io_data_in[7:0] ? 8'h2d : _GEN_505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_507 = 8'hfb == io_data_in[7:0] ? 8'hf : _GEN_506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_508 = 8'hfc == io_data_in[7:0] ? 8'hb0 : _GEN_507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_509 = 8'hfd == io_data_in[7:0] ? 8'h54 : _GEN_508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_510 = 8'hfe == io_data_in[7:0] ? 8'hbb : _GEN_509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_511 = 8'hff == io_data_in[7:0] ? 8'h16 : _GEN_510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_513 = 8'h1 == io_data_in[31:24] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_514 = 8'h2 == io_data_in[31:24] ? 8'h77 : _GEN_513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_515 = 8'h3 == io_data_in[31:24] ? 8'h7b : _GEN_514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_516 = 8'h4 == io_data_in[31:24] ? 8'hf2 : _GEN_515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_517 = 8'h5 == io_data_in[31:24] ? 8'h6b : _GEN_516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_518 = 8'h6 == io_data_in[31:24] ? 8'h6f : _GEN_517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_519 = 8'h7 == io_data_in[31:24] ? 8'hc5 : _GEN_518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_520 = 8'h8 == io_data_in[31:24] ? 8'h30 : _GEN_519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_521 = 8'h9 == io_data_in[31:24] ? 8'h1 : _GEN_520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_522 = 8'ha == io_data_in[31:24] ? 8'h67 : _GEN_521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_523 = 8'hb == io_data_in[31:24] ? 8'h2b : _GEN_522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_524 = 8'hc == io_data_in[31:24] ? 8'hfe : _GEN_523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_525 = 8'hd == io_data_in[31:24] ? 8'hd7 : _GEN_524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_526 = 8'he == io_data_in[31:24] ? 8'hab : _GEN_525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_527 = 8'hf == io_data_in[31:24] ? 8'h76 : _GEN_526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_528 = 8'h10 == io_data_in[31:24] ? 8'hca : _GEN_527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_529 = 8'h11 == io_data_in[31:24] ? 8'h82 : _GEN_528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_530 = 8'h12 == io_data_in[31:24] ? 8'hc9 : _GEN_529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_531 = 8'h13 == io_data_in[31:24] ? 8'h7d : _GEN_530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_532 = 8'h14 == io_data_in[31:24] ? 8'hfa : _GEN_531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_533 = 8'h15 == io_data_in[31:24] ? 8'h59 : _GEN_532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_534 = 8'h16 == io_data_in[31:24] ? 8'h47 : _GEN_533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_535 = 8'h17 == io_data_in[31:24] ? 8'hf0 : _GEN_534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_536 = 8'h18 == io_data_in[31:24] ? 8'had : _GEN_535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_537 = 8'h19 == io_data_in[31:24] ? 8'hd4 : _GEN_536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_538 = 8'h1a == io_data_in[31:24] ? 8'ha2 : _GEN_537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_539 = 8'h1b == io_data_in[31:24] ? 8'haf : _GEN_538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_540 = 8'h1c == io_data_in[31:24] ? 8'h9c : _GEN_539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_541 = 8'h1d == io_data_in[31:24] ? 8'ha4 : _GEN_540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_542 = 8'h1e == io_data_in[31:24] ? 8'h72 : _GEN_541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_543 = 8'h1f == io_data_in[31:24] ? 8'hc0 : _GEN_542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_544 = 8'h20 == io_data_in[31:24] ? 8'hb7 : _GEN_543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_545 = 8'h21 == io_data_in[31:24] ? 8'hfd : _GEN_544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_546 = 8'h22 == io_data_in[31:24] ? 8'h93 : _GEN_545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_547 = 8'h23 == io_data_in[31:24] ? 8'h26 : _GEN_546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_548 = 8'h24 == io_data_in[31:24] ? 8'h36 : _GEN_547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_549 = 8'h25 == io_data_in[31:24] ? 8'h3f : _GEN_548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_550 = 8'h26 == io_data_in[31:24] ? 8'hf7 : _GEN_549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_551 = 8'h27 == io_data_in[31:24] ? 8'hcc : _GEN_550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_552 = 8'h28 == io_data_in[31:24] ? 8'h34 : _GEN_551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_553 = 8'h29 == io_data_in[31:24] ? 8'ha5 : _GEN_552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_554 = 8'h2a == io_data_in[31:24] ? 8'he5 : _GEN_553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_555 = 8'h2b == io_data_in[31:24] ? 8'hf1 : _GEN_554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_556 = 8'h2c == io_data_in[31:24] ? 8'h71 : _GEN_555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_557 = 8'h2d == io_data_in[31:24] ? 8'hd8 : _GEN_556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_558 = 8'h2e == io_data_in[31:24] ? 8'h31 : _GEN_557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_559 = 8'h2f == io_data_in[31:24] ? 8'h15 : _GEN_558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_560 = 8'h30 == io_data_in[31:24] ? 8'h4 : _GEN_559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_561 = 8'h31 == io_data_in[31:24] ? 8'hc7 : _GEN_560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_562 = 8'h32 == io_data_in[31:24] ? 8'h23 : _GEN_561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_563 = 8'h33 == io_data_in[31:24] ? 8'hc3 : _GEN_562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_564 = 8'h34 == io_data_in[31:24] ? 8'h18 : _GEN_563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_565 = 8'h35 == io_data_in[31:24] ? 8'h96 : _GEN_564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_566 = 8'h36 == io_data_in[31:24] ? 8'h5 : _GEN_565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_567 = 8'h37 == io_data_in[31:24] ? 8'h9a : _GEN_566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_568 = 8'h38 == io_data_in[31:24] ? 8'h7 : _GEN_567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_569 = 8'h39 == io_data_in[31:24] ? 8'h12 : _GEN_568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_570 = 8'h3a == io_data_in[31:24] ? 8'h80 : _GEN_569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_571 = 8'h3b == io_data_in[31:24] ? 8'he2 : _GEN_570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_572 = 8'h3c == io_data_in[31:24] ? 8'heb : _GEN_571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_573 = 8'h3d == io_data_in[31:24] ? 8'h27 : _GEN_572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_574 = 8'h3e == io_data_in[31:24] ? 8'hb2 : _GEN_573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_575 = 8'h3f == io_data_in[31:24] ? 8'h75 : _GEN_574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_576 = 8'h40 == io_data_in[31:24] ? 8'h9 : _GEN_575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_577 = 8'h41 == io_data_in[31:24] ? 8'h83 : _GEN_576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_578 = 8'h42 == io_data_in[31:24] ? 8'h2c : _GEN_577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_579 = 8'h43 == io_data_in[31:24] ? 8'h1a : _GEN_578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_580 = 8'h44 == io_data_in[31:24] ? 8'h1b : _GEN_579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_581 = 8'h45 == io_data_in[31:24] ? 8'h6e : _GEN_580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_582 = 8'h46 == io_data_in[31:24] ? 8'h5a : _GEN_581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_583 = 8'h47 == io_data_in[31:24] ? 8'ha0 : _GEN_582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_584 = 8'h48 == io_data_in[31:24] ? 8'h52 : _GEN_583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_585 = 8'h49 == io_data_in[31:24] ? 8'h3b : _GEN_584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_586 = 8'h4a == io_data_in[31:24] ? 8'hd6 : _GEN_585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_587 = 8'h4b == io_data_in[31:24] ? 8'hb3 : _GEN_586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_588 = 8'h4c == io_data_in[31:24] ? 8'h29 : _GEN_587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_589 = 8'h4d == io_data_in[31:24] ? 8'he3 : _GEN_588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_590 = 8'h4e == io_data_in[31:24] ? 8'h2f : _GEN_589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_591 = 8'h4f == io_data_in[31:24] ? 8'h84 : _GEN_590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_592 = 8'h50 == io_data_in[31:24] ? 8'h53 : _GEN_591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_593 = 8'h51 == io_data_in[31:24] ? 8'hd1 : _GEN_592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_594 = 8'h52 == io_data_in[31:24] ? 8'h0 : _GEN_593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_595 = 8'h53 == io_data_in[31:24] ? 8'hed : _GEN_594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_596 = 8'h54 == io_data_in[31:24] ? 8'h20 : _GEN_595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_597 = 8'h55 == io_data_in[31:24] ? 8'hfc : _GEN_596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_598 = 8'h56 == io_data_in[31:24] ? 8'hb1 : _GEN_597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_599 = 8'h57 == io_data_in[31:24] ? 8'h5b : _GEN_598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_600 = 8'h58 == io_data_in[31:24] ? 8'h6a : _GEN_599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_601 = 8'h59 == io_data_in[31:24] ? 8'hcb : _GEN_600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_602 = 8'h5a == io_data_in[31:24] ? 8'hbe : _GEN_601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_603 = 8'h5b == io_data_in[31:24] ? 8'h39 : _GEN_602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_604 = 8'h5c == io_data_in[31:24] ? 8'h4a : _GEN_603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_605 = 8'h5d == io_data_in[31:24] ? 8'h4c : _GEN_604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_606 = 8'h5e == io_data_in[31:24] ? 8'h58 : _GEN_605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_607 = 8'h5f == io_data_in[31:24] ? 8'hcf : _GEN_606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_608 = 8'h60 == io_data_in[31:24] ? 8'hd0 : _GEN_607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_609 = 8'h61 == io_data_in[31:24] ? 8'hef : _GEN_608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_610 = 8'h62 == io_data_in[31:24] ? 8'haa : _GEN_609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_611 = 8'h63 == io_data_in[31:24] ? 8'hfb : _GEN_610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_612 = 8'h64 == io_data_in[31:24] ? 8'h43 : _GEN_611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_613 = 8'h65 == io_data_in[31:24] ? 8'h4d : _GEN_612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_614 = 8'h66 == io_data_in[31:24] ? 8'h33 : _GEN_613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_615 = 8'h67 == io_data_in[31:24] ? 8'h85 : _GEN_614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_616 = 8'h68 == io_data_in[31:24] ? 8'h45 : _GEN_615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_617 = 8'h69 == io_data_in[31:24] ? 8'hf9 : _GEN_616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_618 = 8'h6a == io_data_in[31:24] ? 8'h2 : _GEN_617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_619 = 8'h6b == io_data_in[31:24] ? 8'h7f : _GEN_618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_620 = 8'h6c == io_data_in[31:24] ? 8'h50 : _GEN_619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_621 = 8'h6d == io_data_in[31:24] ? 8'h3c : _GEN_620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_622 = 8'h6e == io_data_in[31:24] ? 8'h9f : _GEN_621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_623 = 8'h6f == io_data_in[31:24] ? 8'ha8 : _GEN_622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_624 = 8'h70 == io_data_in[31:24] ? 8'h51 : _GEN_623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_625 = 8'h71 == io_data_in[31:24] ? 8'ha3 : _GEN_624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_626 = 8'h72 == io_data_in[31:24] ? 8'h40 : _GEN_625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_627 = 8'h73 == io_data_in[31:24] ? 8'h8f : _GEN_626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_628 = 8'h74 == io_data_in[31:24] ? 8'h92 : _GEN_627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_629 = 8'h75 == io_data_in[31:24] ? 8'h9d : _GEN_628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_630 = 8'h76 == io_data_in[31:24] ? 8'h38 : _GEN_629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_631 = 8'h77 == io_data_in[31:24] ? 8'hf5 : _GEN_630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_632 = 8'h78 == io_data_in[31:24] ? 8'hbc : _GEN_631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_633 = 8'h79 == io_data_in[31:24] ? 8'hb6 : _GEN_632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_634 = 8'h7a == io_data_in[31:24] ? 8'hda : _GEN_633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_635 = 8'h7b == io_data_in[31:24] ? 8'h21 : _GEN_634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_636 = 8'h7c == io_data_in[31:24] ? 8'h10 : _GEN_635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_637 = 8'h7d == io_data_in[31:24] ? 8'hff : _GEN_636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_638 = 8'h7e == io_data_in[31:24] ? 8'hf3 : _GEN_637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_639 = 8'h7f == io_data_in[31:24] ? 8'hd2 : _GEN_638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_640 = 8'h80 == io_data_in[31:24] ? 8'hcd : _GEN_639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_641 = 8'h81 == io_data_in[31:24] ? 8'hc : _GEN_640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_642 = 8'h82 == io_data_in[31:24] ? 8'h13 : _GEN_641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_643 = 8'h83 == io_data_in[31:24] ? 8'hec : _GEN_642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_644 = 8'h84 == io_data_in[31:24] ? 8'h5f : _GEN_643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_645 = 8'h85 == io_data_in[31:24] ? 8'h97 : _GEN_644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_646 = 8'h86 == io_data_in[31:24] ? 8'h44 : _GEN_645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_647 = 8'h87 == io_data_in[31:24] ? 8'h17 : _GEN_646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_648 = 8'h88 == io_data_in[31:24] ? 8'hc4 : _GEN_647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_649 = 8'h89 == io_data_in[31:24] ? 8'ha7 : _GEN_648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_650 = 8'h8a == io_data_in[31:24] ? 8'h7e : _GEN_649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_651 = 8'h8b == io_data_in[31:24] ? 8'h3d : _GEN_650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_652 = 8'h8c == io_data_in[31:24] ? 8'h64 : _GEN_651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_653 = 8'h8d == io_data_in[31:24] ? 8'h5d : _GEN_652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_654 = 8'h8e == io_data_in[31:24] ? 8'h19 : _GEN_653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_655 = 8'h8f == io_data_in[31:24] ? 8'h73 : _GEN_654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_656 = 8'h90 == io_data_in[31:24] ? 8'h60 : _GEN_655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_657 = 8'h91 == io_data_in[31:24] ? 8'h81 : _GEN_656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_658 = 8'h92 == io_data_in[31:24] ? 8'h4f : _GEN_657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_659 = 8'h93 == io_data_in[31:24] ? 8'hdc : _GEN_658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_660 = 8'h94 == io_data_in[31:24] ? 8'h22 : _GEN_659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_661 = 8'h95 == io_data_in[31:24] ? 8'h2a : _GEN_660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_662 = 8'h96 == io_data_in[31:24] ? 8'h90 : _GEN_661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_663 = 8'h97 == io_data_in[31:24] ? 8'h88 : _GEN_662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_664 = 8'h98 == io_data_in[31:24] ? 8'h46 : _GEN_663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_665 = 8'h99 == io_data_in[31:24] ? 8'hee : _GEN_664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_666 = 8'h9a == io_data_in[31:24] ? 8'hb8 : _GEN_665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_667 = 8'h9b == io_data_in[31:24] ? 8'h14 : _GEN_666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_668 = 8'h9c == io_data_in[31:24] ? 8'hde : _GEN_667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_669 = 8'h9d == io_data_in[31:24] ? 8'h5e : _GEN_668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_670 = 8'h9e == io_data_in[31:24] ? 8'hb : _GEN_669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_671 = 8'h9f == io_data_in[31:24] ? 8'hdb : _GEN_670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_672 = 8'ha0 == io_data_in[31:24] ? 8'he0 : _GEN_671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_673 = 8'ha1 == io_data_in[31:24] ? 8'h32 : _GEN_672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_674 = 8'ha2 == io_data_in[31:24] ? 8'h3a : _GEN_673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_675 = 8'ha3 == io_data_in[31:24] ? 8'ha : _GEN_674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_676 = 8'ha4 == io_data_in[31:24] ? 8'h49 : _GEN_675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_677 = 8'ha5 == io_data_in[31:24] ? 8'h6 : _GEN_676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_678 = 8'ha6 == io_data_in[31:24] ? 8'h24 : _GEN_677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_679 = 8'ha7 == io_data_in[31:24] ? 8'h5c : _GEN_678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_680 = 8'ha8 == io_data_in[31:24] ? 8'hc2 : _GEN_679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_681 = 8'ha9 == io_data_in[31:24] ? 8'hd3 : _GEN_680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_682 = 8'haa == io_data_in[31:24] ? 8'hac : _GEN_681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_683 = 8'hab == io_data_in[31:24] ? 8'h62 : _GEN_682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_684 = 8'hac == io_data_in[31:24] ? 8'h91 : _GEN_683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_685 = 8'had == io_data_in[31:24] ? 8'h95 : _GEN_684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_686 = 8'hae == io_data_in[31:24] ? 8'he4 : _GEN_685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_687 = 8'haf == io_data_in[31:24] ? 8'h79 : _GEN_686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_688 = 8'hb0 == io_data_in[31:24] ? 8'he7 : _GEN_687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_689 = 8'hb1 == io_data_in[31:24] ? 8'hc8 : _GEN_688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_690 = 8'hb2 == io_data_in[31:24] ? 8'h37 : _GEN_689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_691 = 8'hb3 == io_data_in[31:24] ? 8'h6d : _GEN_690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_692 = 8'hb4 == io_data_in[31:24] ? 8'h8d : _GEN_691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_693 = 8'hb5 == io_data_in[31:24] ? 8'hd5 : _GEN_692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_694 = 8'hb6 == io_data_in[31:24] ? 8'h4e : _GEN_693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_695 = 8'hb7 == io_data_in[31:24] ? 8'ha9 : _GEN_694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_696 = 8'hb8 == io_data_in[31:24] ? 8'h6c : _GEN_695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_697 = 8'hb9 == io_data_in[31:24] ? 8'h56 : _GEN_696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_698 = 8'hba == io_data_in[31:24] ? 8'hf4 : _GEN_697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_699 = 8'hbb == io_data_in[31:24] ? 8'hea : _GEN_698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_700 = 8'hbc == io_data_in[31:24] ? 8'h65 : _GEN_699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_701 = 8'hbd == io_data_in[31:24] ? 8'h7a : _GEN_700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_702 = 8'hbe == io_data_in[31:24] ? 8'hae : _GEN_701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_703 = 8'hbf == io_data_in[31:24] ? 8'h8 : _GEN_702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_704 = 8'hc0 == io_data_in[31:24] ? 8'hba : _GEN_703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_705 = 8'hc1 == io_data_in[31:24] ? 8'h78 : _GEN_704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_706 = 8'hc2 == io_data_in[31:24] ? 8'h25 : _GEN_705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_707 = 8'hc3 == io_data_in[31:24] ? 8'h2e : _GEN_706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_708 = 8'hc4 == io_data_in[31:24] ? 8'h1c : _GEN_707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_709 = 8'hc5 == io_data_in[31:24] ? 8'ha6 : _GEN_708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_710 = 8'hc6 == io_data_in[31:24] ? 8'hb4 : _GEN_709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_711 = 8'hc7 == io_data_in[31:24] ? 8'hc6 : _GEN_710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_712 = 8'hc8 == io_data_in[31:24] ? 8'he8 : _GEN_711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_713 = 8'hc9 == io_data_in[31:24] ? 8'hdd : _GEN_712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_714 = 8'hca == io_data_in[31:24] ? 8'h74 : _GEN_713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_715 = 8'hcb == io_data_in[31:24] ? 8'h1f : _GEN_714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_716 = 8'hcc == io_data_in[31:24] ? 8'h4b : _GEN_715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_717 = 8'hcd == io_data_in[31:24] ? 8'hbd : _GEN_716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_718 = 8'hce == io_data_in[31:24] ? 8'h8b : _GEN_717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_719 = 8'hcf == io_data_in[31:24] ? 8'h8a : _GEN_718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_720 = 8'hd0 == io_data_in[31:24] ? 8'h70 : _GEN_719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_721 = 8'hd1 == io_data_in[31:24] ? 8'h3e : _GEN_720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_722 = 8'hd2 == io_data_in[31:24] ? 8'hb5 : _GEN_721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_723 = 8'hd3 == io_data_in[31:24] ? 8'h66 : _GEN_722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_724 = 8'hd4 == io_data_in[31:24] ? 8'h48 : _GEN_723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_725 = 8'hd5 == io_data_in[31:24] ? 8'h3 : _GEN_724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_726 = 8'hd6 == io_data_in[31:24] ? 8'hf6 : _GEN_725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_727 = 8'hd7 == io_data_in[31:24] ? 8'he : _GEN_726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_728 = 8'hd8 == io_data_in[31:24] ? 8'h61 : _GEN_727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_729 = 8'hd9 == io_data_in[31:24] ? 8'h35 : _GEN_728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_730 = 8'hda == io_data_in[31:24] ? 8'h57 : _GEN_729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_731 = 8'hdb == io_data_in[31:24] ? 8'hb9 : _GEN_730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_732 = 8'hdc == io_data_in[31:24] ? 8'h86 : _GEN_731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_733 = 8'hdd == io_data_in[31:24] ? 8'hc1 : _GEN_732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_734 = 8'hde == io_data_in[31:24] ? 8'h1d : _GEN_733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_735 = 8'hdf == io_data_in[31:24] ? 8'h9e : _GEN_734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_736 = 8'he0 == io_data_in[31:24] ? 8'he1 : _GEN_735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_737 = 8'he1 == io_data_in[31:24] ? 8'hf8 : _GEN_736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_738 = 8'he2 == io_data_in[31:24] ? 8'h98 : _GEN_737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_739 = 8'he3 == io_data_in[31:24] ? 8'h11 : _GEN_738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_740 = 8'he4 == io_data_in[31:24] ? 8'h69 : _GEN_739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_741 = 8'he5 == io_data_in[31:24] ? 8'hd9 : _GEN_740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_742 = 8'he6 == io_data_in[31:24] ? 8'h8e : _GEN_741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_743 = 8'he7 == io_data_in[31:24] ? 8'h94 : _GEN_742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_744 = 8'he8 == io_data_in[31:24] ? 8'h9b : _GEN_743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_745 = 8'he9 == io_data_in[31:24] ? 8'h1e : _GEN_744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_746 = 8'hea == io_data_in[31:24] ? 8'h87 : _GEN_745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_747 = 8'heb == io_data_in[31:24] ? 8'he9 : _GEN_746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_748 = 8'hec == io_data_in[31:24] ? 8'hce : _GEN_747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_749 = 8'hed == io_data_in[31:24] ? 8'h55 : _GEN_748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_750 = 8'hee == io_data_in[31:24] ? 8'h28 : _GEN_749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_751 = 8'hef == io_data_in[31:24] ? 8'hdf : _GEN_750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_752 = 8'hf0 == io_data_in[31:24] ? 8'h8c : _GEN_751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_753 = 8'hf1 == io_data_in[31:24] ? 8'ha1 : _GEN_752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_754 = 8'hf2 == io_data_in[31:24] ? 8'h89 : _GEN_753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_755 = 8'hf3 == io_data_in[31:24] ? 8'hd : _GEN_754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_756 = 8'hf4 == io_data_in[31:24] ? 8'hbf : _GEN_755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_757 = 8'hf5 == io_data_in[31:24] ? 8'he6 : _GEN_756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_758 = 8'hf6 == io_data_in[31:24] ? 8'h42 : _GEN_757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_759 = 8'hf7 == io_data_in[31:24] ? 8'h68 : _GEN_758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_760 = 8'hf8 == io_data_in[31:24] ? 8'h41 : _GEN_759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_761 = 8'hf9 == io_data_in[31:24] ? 8'h99 : _GEN_760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_762 = 8'hfa == io_data_in[31:24] ? 8'h2d : _GEN_761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_763 = 8'hfb == io_data_in[31:24] ? 8'hf : _GEN_762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_764 = 8'hfc == io_data_in[31:24] ? 8'hb0 : _GEN_763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_765 = 8'hfd == io_data_in[31:24] ? 8'h54 : _GEN_764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_766 = 8'hfe == io_data_in[31:24] ? 8'hbb : _GEN_765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_767 = 8'hff == io_data_in[31:24] ? 8'h16 : _GEN_766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_769 = 8'h1 == io_data_in[23:16] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_770 = 8'h2 == io_data_in[23:16] ? 8'h77 : _GEN_769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_771 = 8'h3 == io_data_in[23:16] ? 8'h7b : _GEN_770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_772 = 8'h4 == io_data_in[23:16] ? 8'hf2 : _GEN_771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_773 = 8'h5 == io_data_in[23:16] ? 8'h6b : _GEN_772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_774 = 8'h6 == io_data_in[23:16] ? 8'h6f : _GEN_773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_775 = 8'h7 == io_data_in[23:16] ? 8'hc5 : _GEN_774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_776 = 8'h8 == io_data_in[23:16] ? 8'h30 : _GEN_775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_777 = 8'h9 == io_data_in[23:16] ? 8'h1 : _GEN_776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_778 = 8'ha == io_data_in[23:16] ? 8'h67 : _GEN_777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_779 = 8'hb == io_data_in[23:16] ? 8'h2b : _GEN_778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_780 = 8'hc == io_data_in[23:16] ? 8'hfe : _GEN_779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_781 = 8'hd == io_data_in[23:16] ? 8'hd7 : _GEN_780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_782 = 8'he == io_data_in[23:16] ? 8'hab : _GEN_781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_783 = 8'hf == io_data_in[23:16] ? 8'h76 : _GEN_782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_784 = 8'h10 == io_data_in[23:16] ? 8'hca : _GEN_783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_785 = 8'h11 == io_data_in[23:16] ? 8'h82 : _GEN_784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_786 = 8'h12 == io_data_in[23:16] ? 8'hc9 : _GEN_785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_787 = 8'h13 == io_data_in[23:16] ? 8'h7d : _GEN_786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_788 = 8'h14 == io_data_in[23:16] ? 8'hfa : _GEN_787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_789 = 8'h15 == io_data_in[23:16] ? 8'h59 : _GEN_788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_790 = 8'h16 == io_data_in[23:16] ? 8'h47 : _GEN_789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_791 = 8'h17 == io_data_in[23:16] ? 8'hf0 : _GEN_790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_792 = 8'h18 == io_data_in[23:16] ? 8'had : _GEN_791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_793 = 8'h19 == io_data_in[23:16] ? 8'hd4 : _GEN_792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_794 = 8'h1a == io_data_in[23:16] ? 8'ha2 : _GEN_793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_795 = 8'h1b == io_data_in[23:16] ? 8'haf : _GEN_794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_796 = 8'h1c == io_data_in[23:16] ? 8'h9c : _GEN_795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_797 = 8'h1d == io_data_in[23:16] ? 8'ha4 : _GEN_796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_798 = 8'h1e == io_data_in[23:16] ? 8'h72 : _GEN_797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_799 = 8'h1f == io_data_in[23:16] ? 8'hc0 : _GEN_798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_800 = 8'h20 == io_data_in[23:16] ? 8'hb7 : _GEN_799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_801 = 8'h21 == io_data_in[23:16] ? 8'hfd : _GEN_800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_802 = 8'h22 == io_data_in[23:16] ? 8'h93 : _GEN_801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_803 = 8'h23 == io_data_in[23:16] ? 8'h26 : _GEN_802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_804 = 8'h24 == io_data_in[23:16] ? 8'h36 : _GEN_803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_805 = 8'h25 == io_data_in[23:16] ? 8'h3f : _GEN_804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_806 = 8'h26 == io_data_in[23:16] ? 8'hf7 : _GEN_805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_807 = 8'h27 == io_data_in[23:16] ? 8'hcc : _GEN_806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_808 = 8'h28 == io_data_in[23:16] ? 8'h34 : _GEN_807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_809 = 8'h29 == io_data_in[23:16] ? 8'ha5 : _GEN_808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_810 = 8'h2a == io_data_in[23:16] ? 8'he5 : _GEN_809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_811 = 8'h2b == io_data_in[23:16] ? 8'hf1 : _GEN_810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_812 = 8'h2c == io_data_in[23:16] ? 8'h71 : _GEN_811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_813 = 8'h2d == io_data_in[23:16] ? 8'hd8 : _GEN_812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_814 = 8'h2e == io_data_in[23:16] ? 8'h31 : _GEN_813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_815 = 8'h2f == io_data_in[23:16] ? 8'h15 : _GEN_814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_816 = 8'h30 == io_data_in[23:16] ? 8'h4 : _GEN_815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_817 = 8'h31 == io_data_in[23:16] ? 8'hc7 : _GEN_816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_818 = 8'h32 == io_data_in[23:16] ? 8'h23 : _GEN_817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_819 = 8'h33 == io_data_in[23:16] ? 8'hc3 : _GEN_818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_820 = 8'h34 == io_data_in[23:16] ? 8'h18 : _GEN_819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_821 = 8'h35 == io_data_in[23:16] ? 8'h96 : _GEN_820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_822 = 8'h36 == io_data_in[23:16] ? 8'h5 : _GEN_821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_823 = 8'h37 == io_data_in[23:16] ? 8'h9a : _GEN_822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_824 = 8'h38 == io_data_in[23:16] ? 8'h7 : _GEN_823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_825 = 8'h39 == io_data_in[23:16] ? 8'h12 : _GEN_824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_826 = 8'h3a == io_data_in[23:16] ? 8'h80 : _GEN_825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_827 = 8'h3b == io_data_in[23:16] ? 8'he2 : _GEN_826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_828 = 8'h3c == io_data_in[23:16] ? 8'heb : _GEN_827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_829 = 8'h3d == io_data_in[23:16] ? 8'h27 : _GEN_828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_830 = 8'h3e == io_data_in[23:16] ? 8'hb2 : _GEN_829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_831 = 8'h3f == io_data_in[23:16] ? 8'h75 : _GEN_830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_832 = 8'h40 == io_data_in[23:16] ? 8'h9 : _GEN_831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_833 = 8'h41 == io_data_in[23:16] ? 8'h83 : _GEN_832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_834 = 8'h42 == io_data_in[23:16] ? 8'h2c : _GEN_833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_835 = 8'h43 == io_data_in[23:16] ? 8'h1a : _GEN_834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_836 = 8'h44 == io_data_in[23:16] ? 8'h1b : _GEN_835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_837 = 8'h45 == io_data_in[23:16] ? 8'h6e : _GEN_836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_838 = 8'h46 == io_data_in[23:16] ? 8'h5a : _GEN_837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_839 = 8'h47 == io_data_in[23:16] ? 8'ha0 : _GEN_838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_840 = 8'h48 == io_data_in[23:16] ? 8'h52 : _GEN_839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_841 = 8'h49 == io_data_in[23:16] ? 8'h3b : _GEN_840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_842 = 8'h4a == io_data_in[23:16] ? 8'hd6 : _GEN_841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_843 = 8'h4b == io_data_in[23:16] ? 8'hb3 : _GEN_842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_844 = 8'h4c == io_data_in[23:16] ? 8'h29 : _GEN_843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_845 = 8'h4d == io_data_in[23:16] ? 8'he3 : _GEN_844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_846 = 8'h4e == io_data_in[23:16] ? 8'h2f : _GEN_845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_847 = 8'h4f == io_data_in[23:16] ? 8'h84 : _GEN_846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_848 = 8'h50 == io_data_in[23:16] ? 8'h53 : _GEN_847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_849 = 8'h51 == io_data_in[23:16] ? 8'hd1 : _GEN_848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_850 = 8'h52 == io_data_in[23:16] ? 8'h0 : _GEN_849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_851 = 8'h53 == io_data_in[23:16] ? 8'hed : _GEN_850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_852 = 8'h54 == io_data_in[23:16] ? 8'h20 : _GEN_851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_853 = 8'h55 == io_data_in[23:16] ? 8'hfc : _GEN_852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_854 = 8'h56 == io_data_in[23:16] ? 8'hb1 : _GEN_853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_855 = 8'h57 == io_data_in[23:16] ? 8'h5b : _GEN_854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_856 = 8'h58 == io_data_in[23:16] ? 8'h6a : _GEN_855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_857 = 8'h59 == io_data_in[23:16] ? 8'hcb : _GEN_856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_858 = 8'h5a == io_data_in[23:16] ? 8'hbe : _GEN_857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_859 = 8'h5b == io_data_in[23:16] ? 8'h39 : _GEN_858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_860 = 8'h5c == io_data_in[23:16] ? 8'h4a : _GEN_859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_861 = 8'h5d == io_data_in[23:16] ? 8'h4c : _GEN_860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_862 = 8'h5e == io_data_in[23:16] ? 8'h58 : _GEN_861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_863 = 8'h5f == io_data_in[23:16] ? 8'hcf : _GEN_862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_864 = 8'h60 == io_data_in[23:16] ? 8'hd0 : _GEN_863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_865 = 8'h61 == io_data_in[23:16] ? 8'hef : _GEN_864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_866 = 8'h62 == io_data_in[23:16] ? 8'haa : _GEN_865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_867 = 8'h63 == io_data_in[23:16] ? 8'hfb : _GEN_866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_868 = 8'h64 == io_data_in[23:16] ? 8'h43 : _GEN_867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_869 = 8'h65 == io_data_in[23:16] ? 8'h4d : _GEN_868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_870 = 8'h66 == io_data_in[23:16] ? 8'h33 : _GEN_869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_871 = 8'h67 == io_data_in[23:16] ? 8'h85 : _GEN_870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_872 = 8'h68 == io_data_in[23:16] ? 8'h45 : _GEN_871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_873 = 8'h69 == io_data_in[23:16] ? 8'hf9 : _GEN_872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_874 = 8'h6a == io_data_in[23:16] ? 8'h2 : _GEN_873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_875 = 8'h6b == io_data_in[23:16] ? 8'h7f : _GEN_874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_876 = 8'h6c == io_data_in[23:16] ? 8'h50 : _GEN_875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_877 = 8'h6d == io_data_in[23:16] ? 8'h3c : _GEN_876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_878 = 8'h6e == io_data_in[23:16] ? 8'h9f : _GEN_877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_879 = 8'h6f == io_data_in[23:16] ? 8'ha8 : _GEN_878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_880 = 8'h70 == io_data_in[23:16] ? 8'h51 : _GEN_879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_881 = 8'h71 == io_data_in[23:16] ? 8'ha3 : _GEN_880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_882 = 8'h72 == io_data_in[23:16] ? 8'h40 : _GEN_881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_883 = 8'h73 == io_data_in[23:16] ? 8'h8f : _GEN_882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_884 = 8'h74 == io_data_in[23:16] ? 8'h92 : _GEN_883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_885 = 8'h75 == io_data_in[23:16] ? 8'h9d : _GEN_884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_886 = 8'h76 == io_data_in[23:16] ? 8'h38 : _GEN_885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_887 = 8'h77 == io_data_in[23:16] ? 8'hf5 : _GEN_886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_888 = 8'h78 == io_data_in[23:16] ? 8'hbc : _GEN_887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_889 = 8'h79 == io_data_in[23:16] ? 8'hb6 : _GEN_888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_890 = 8'h7a == io_data_in[23:16] ? 8'hda : _GEN_889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_891 = 8'h7b == io_data_in[23:16] ? 8'h21 : _GEN_890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_892 = 8'h7c == io_data_in[23:16] ? 8'h10 : _GEN_891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_893 = 8'h7d == io_data_in[23:16] ? 8'hff : _GEN_892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_894 = 8'h7e == io_data_in[23:16] ? 8'hf3 : _GEN_893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_895 = 8'h7f == io_data_in[23:16] ? 8'hd2 : _GEN_894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_896 = 8'h80 == io_data_in[23:16] ? 8'hcd : _GEN_895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_897 = 8'h81 == io_data_in[23:16] ? 8'hc : _GEN_896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_898 = 8'h82 == io_data_in[23:16] ? 8'h13 : _GEN_897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_899 = 8'h83 == io_data_in[23:16] ? 8'hec : _GEN_898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_900 = 8'h84 == io_data_in[23:16] ? 8'h5f : _GEN_899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_901 = 8'h85 == io_data_in[23:16] ? 8'h97 : _GEN_900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_902 = 8'h86 == io_data_in[23:16] ? 8'h44 : _GEN_901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_903 = 8'h87 == io_data_in[23:16] ? 8'h17 : _GEN_902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_904 = 8'h88 == io_data_in[23:16] ? 8'hc4 : _GEN_903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_905 = 8'h89 == io_data_in[23:16] ? 8'ha7 : _GEN_904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_906 = 8'h8a == io_data_in[23:16] ? 8'h7e : _GEN_905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_907 = 8'h8b == io_data_in[23:16] ? 8'h3d : _GEN_906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_908 = 8'h8c == io_data_in[23:16] ? 8'h64 : _GEN_907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_909 = 8'h8d == io_data_in[23:16] ? 8'h5d : _GEN_908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_910 = 8'h8e == io_data_in[23:16] ? 8'h19 : _GEN_909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_911 = 8'h8f == io_data_in[23:16] ? 8'h73 : _GEN_910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_912 = 8'h90 == io_data_in[23:16] ? 8'h60 : _GEN_911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_913 = 8'h91 == io_data_in[23:16] ? 8'h81 : _GEN_912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_914 = 8'h92 == io_data_in[23:16] ? 8'h4f : _GEN_913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_915 = 8'h93 == io_data_in[23:16] ? 8'hdc : _GEN_914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_916 = 8'h94 == io_data_in[23:16] ? 8'h22 : _GEN_915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_917 = 8'h95 == io_data_in[23:16] ? 8'h2a : _GEN_916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_918 = 8'h96 == io_data_in[23:16] ? 8'h90 : _GEN_917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_919 = 8'h97 == io_data_in[23:16] ? 8'h88 : _GEN_918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_920 = 8'h98 == io_data_in[23:16] ? 8'h46 : _GEN_919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_921 = 8'h99 == io_data_in[23:16] ? 8'hee : _GEN_920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_922 = 8'h9a == io_data_in[23:16] ? 8'hb8 : _GEN_921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_923 = 8'h9b == io_data_in[23:16] ? 8'h14 : _GEN_922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_924 = 8'h9c == io_data_in[23:16] ? 8'hde : _GEN_923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_925 = 8'h9d == io_data_in[23:16] ? 8'h5e : _GEN_924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_926 = 8'h9e == io_data_in[23:16] ? 8'hb : _GEN_925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_927 = 8'h9f == io_data_in[23:16] ? 8'hdb : _GEN_926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_928 = 8'ha0 == io_data_in[23:16] ? 8'he0 : _GEN_927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_929 = 8'ha1 == io_data_in[23:16] ? 8'h32 : _GEN_928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_930 = 8'ha2 == io_data_in[23:16] ? 8'h3a : _GEN_929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_931 = 8'ha3 == io_data_in[23:16] ? 8'ha : _GEN_930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_932 = 8'ha4 == io_data_in[23:16] ? 8'h49 : _GEN_931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_933 = 8'ha5 == io_data_in[23:16] ? 8'h6 : _GEN_932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_934 = 8'ha6 == io_data_in[23:16] ? 8'h24 : _GEN_933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_935 = 8'ha7 == io_data_in[23:16] ? 8'h5c : _GEN_934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_936 = 8'ha8 == io_data_in[23:16] ? 8'hc2 : _GEN_935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_937 = 8'ha9 == io_data_in[23:16] ? 8'hd3 : _GEN_936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_938 = 8'haa == io_data_in[23:16] ? 8'hac : _GEN_937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_939 = 8'hab == io_data_in[23:16] ? 8'h62 : _GEN_938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_940 = 8'hac == io_data_in[23:16] ? 8'h91 : _GEN_939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_941 = 8'had == io_data_in[23:16] ? 8'h95 : _GEN_940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_942 = 8'hae == io_data_in[23:16] ? 8'he4 : _GEN_941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_943 = 8'haf == io_data_in[23:16] ? 8'h79 : _GEN_942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_944 = 8'hb0 == io_data_in[23:16] ? 8'he7 : _GEN_943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_945 = 8'hb1 == io_data_in[23:16] ? 8'hc8 : _GEN_944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_946 = 8'hb2 == io_data_in[23:16] ? 8'h37 : _GEN_945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_947 = 8'hb3 == io_data_in[23:16] ? 8'h6d : _GEN_946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_948 = 8'hb4 == io_data_in[23:16] ? 8'h8d : _GEN_947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_949 = 8'hb5 == io_data_in[23:16] ? 8'hd5 : _GEN_948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_950 = 8'hb6 == io_data_in[23:16] ? 8'h4e : _GEN_949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_951 = 8'hb7 == io_data_in[23:16] ? 8'ha9 : _GEN_950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_952 = 8'hb8 == io_data_in[23:16] ? 8'h6c : _GEN_951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_953 = 8'hb9 == io_data_in[23:16] ? 8'h56 : _GEN_952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_954 = 8'hba == io_data_in[23:16] ? 8'hf4 : _GEN_953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_955 = 8'hbb == io_data_in[23:16] ? 8'hea : _GEN_954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_956 = 8'hbc == io_data_in[23:16] ? 8'h65 : _GEN_955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_957 = 8'hbd == io_data_in[23:16] ? 8'h7a : _GEN_956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_958 = 8'hbe == io_data_in[23:16] ? 8'hae : _GEN_957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_959 = 8'hbf == io_data_in[23:16] ? 8'h8 : _GEN_958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_960 = 8'hc0 == io_data_in[23:16] ? 8'hba : _GEN_959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_961 = 8'hc1 == io_data_in[23:16] ? 8'h78 : _GEN_960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_962 = 8'hc2 == io_data_in[23:16] ? 8'h25 : _GEN_961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_963 = 8'hc3 == io_data_in[23:16] ? 8'h2e : _GEN_962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_964 = 8'hc4 == io_data_in[23:16] ? 8'h1c : _GEN_963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_965 = 8'hc5 == io_data_in[23:16] ? 8'ha6 : _GEN_964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_966 = 8'hc6 == io_data_in[23:16] ? 8'hb4 : _GEN_965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_967 = 8'hc7 == io_data_in[23:16] ? 8'hc6 : _GEN_966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_968 = 8'hc8 == io_data_in[23:16] ? 8'he8 : _GEN_967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_969 = 8'hc9 == io_data_in[23:16] ? 8'hdd : _GEN_968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_970 = 8'hca == io_data_in[23:16] ? 8'h74 : _GEN_969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_971 = 8'hcb == io_data_in[23:16] ? 8'h1f : _GEN_970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_972 = 8'hcc == io_data_in[23:16] ? 8'h4b : _GEN_971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_973 = 8'hcd == io_data_in[23:16] ? 8'hbd : _GEN_972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_974 = 8'hce == io_data_in[23:16] ? 8'h8b : _GEN_973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_975 = 8'hcf == io_data_in[23:16] ? 8'h8a : _GEN_974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_976 = 8'hd0 == io_data_in[23:16] ? 8'h70 : _GEN_975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_977 = 8'hd1 == io_data_in[23:16] ? 8'h3e : _GEN_976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_978 = 8'hd2 == io_data_in[23:16] ? 8'hb5 : _GEN_977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_979 = 8'hd3 == io_data_in[23:16] ? 8'h66 : _GEN_978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_980 = 8'hd4 == io_data_in[23:16] ? 8'h48 : _GEN_979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_981 = 8'hd5 == io_data_in[23:16] ? 8'h3 : _GEN_980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_982 = 8'hd6 == io_data_in[23:16] ? 8'hf6 : _GEN_981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_983 = 8'hd7 == io_data_in[23:16] ? 8'he : _GEN_982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_984 = 8'hd8 == io_data_in[23:16] ? 8'h61 : _GEN_983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_985 = 8'hd9 == io_data_in[23:16] ? 8'h35 : _GEN_984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_986 = 8'hda == io_data_in[23:16] ? 8'h57 : _GEN_985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_987 = 8'hdb == io_data_in[23:16] ? 8'hb9 : _GEN_986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_988 = 8'hdc == io_data_in[23:16] ? 8'h86 : _GEN_987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_989 = 8'hdd == io_data_in[23:16] ? 8'hc1 : _GEN_988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_990 = 8'hde == io_data_in[23:16] ? 8'h1d : _GEN_989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_991 = 8'hdf == io_data_in[23:16] ? 8'h9e : _GEN_990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_992 = 8'he0 == io_data_in[23:16] ? 8'he1 : _GEN_991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_993 = 8'he1 == io_data_in[23:16] ? 8'hf8 : _GEN_992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_994 = 8'he2 == io_data_in[23:16] ? 8'h98 : _GEN_993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_995 = 8'he3 == io_data_in[23:16] ? 8'h11 : _GEN_994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_996 = 8'he4 == io_data_in[23:16] ? 8'h69 : _GEN_995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_997 = 8'he5 == io_data_in[23:16] ? 8'hd9 : _GEN_996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_998 = 8'he6 == io_data_in[23:16] ? 8'h8e : _GEN_997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_999 = 8'he7 == io_data_in[23:16] ? 8'h94 : _GEN_998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1000 = 8'he8 == io_data_in[23:16] ? 8'h9b : _GEN_999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1001 = 8'he9 == io_data_in[23:16] ? 8'h1e : _GEN_1000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1002 = 8'hea == io_data_in[23:16] ? 8'h87 : _GEN_1001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1003 = 8'heb == io_data_in[23:16] ? 8'he9 : _GEN_1002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1004 = 8'hec == io_data_in[23:16] ? 8'hce : _GEN_1003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1005 = 8'hed == io_data_in[23:16] ? 8'h55 : _GEN_1004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1006 = 8'hee == io_data_in[23:16] ? 8'h28 : _GEN_1005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1007 = 8'hef == io_data_in[23:16] ? 8'hdf : _GEN_1006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1008 = 8'hf0 == io_data_in[23:16] ? 8'h8c : _GEN_1007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1009 = 8'hf1 == io_data_in[23:16] ? 8'ha1 : _GEN_1008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1010 = 8'hf2 == io_data_in[23:16] ? 8'h89 : _GEN_1009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1011 = 8'hf3 == io_data_in[23:16] ? 8'hd : _GEN_1010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1012 = 8'hf4 == io_data_in[23:16] ? 8'hbf : _GEN_1011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1013 = 8'hf5 == io_data_in[23:16] ? 8'he6 : _GEN_1012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1014 = 8'hf6 == io_data_in[23:16] ? 8'h42 : _GEN_1013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1015 = 8'hf7 == io_data_in[23:16] ? 8'h68 : _GEN_1014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1016 = 8'hf8 == io_data_in[23:16] ? 8'h41 : _GEN_1015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1017 = 8'hf9 == io_data_in[23:16] ? 8'h99 : _GEN_1016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1018 = 8'hfa == io_data_in[23:16] ? 8'h2d : _GEN_1017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1019 = 8'hfb == io_data_in[23:16] ? 8'hf : _GEN_1018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1020 = 8'hfc == io_data_in[23:16] ? 8'hb0 : _GEN_1019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1021 = 8'hfd == io_data_in[23:16] ? 8'h54 : _GEN_1020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1022 = 8'hfe == io_data_in[23:16] ? 8'hbb : _GEN_1021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1023 = 8'hff == io_data_in[23:16] ? 8'h16 : _GEN_1022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1025 = 8'h1 == io_data_in[47:40] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1026 = 8'h2 == io_data_in[47:40] ? 8'h77 : _GEN_1025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1027 = 8'h3 == io_data_in[47:40] ? 8'h7b : _GEN_1026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1028 = 8'h4 == io_data_in[47:40] ? 8'hf2 : _GEN_1027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1029 = 8'h5 == io_data_in[47:40] ? 8'h6b : _GEN_1028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1030 = 8'h6 == io_data_in[47:40] ? 8'h6f : _GEN_1029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1031 = 8'h7 == io_data_in[47:40] ? 8'hc5 : _GEN_1030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1032 = 8'h8 == io_data_in[47:40] ? 8'h30 : _GEN_1031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1033 = 8'h9 == io_data_in[47:40] ? 8'h1 : _GEN_1032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1034 = 8'ha == io_data_in[47:40] ? 8'h67 : _GEN_1033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1035 = 8'hb == io_data_in[47:40] ? 8'h2b : _GEN_1034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1036 = 8'hc == io_data_in[47:40] ? 8'hfe : _GEN_1035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1037 = 8'hd == io_data_in[47:40] ? 8'hd7 : _GEN_1036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1038 = 8'he == io_data_in[47:40] ? 8'hab : _GEN_1037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1039 = 8'hf == io_data_in[47:40] ? 8'h76 : _GEN_1038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1040 = 8'h10 == io_data_in[47:40] ? 8'hca : _GEN_1039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1041 = 8'h11 == io_data_in[47:40] ? 8'h82 : _GEN_1040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1042 = 8'h12 == io_data_in[47:40] ? 8'hc9 : _GEN_1041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1043 = 8'h13 == io_data_in[47:40] ? 8'h7d : _GEN_1042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1044 = 8'h14 == io_data_in[47:40] ? 8'hfa : _GEN_1043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1045 = 8'h15 == io_data_in[47:40] ? 8'h59 : _GEN_1044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1046 = 8'h16 == io_data_in[47:40] ? 8'h47 : _GEN_1045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1047 = 8'h17 == io_data_in[47:40] ? 8'hf0 : _GEN_1046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1048 = 8'h18 == io_data_in[47:40] ? 8'had : _GEN_1047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1049 = 8'h19 == io_data_in[47:40] ? 8'hd4 : _GEN_1048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1050 = 8'h1a == io_data_in[47:40] ? 8'ha2 : _GEN_1049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1051 = 8'h1b == io_data_in[47:40] ? 8'haf : _GEN_1050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1052 = 8'h1c == io_data_in[47:40] ? 8'h9c : _GEN_1051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1053 = 8'h1d == io_data_in[47:40] ? 8'ha4 : _GEN_1052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1054 = 8'h1e == io_data_in[47:40] ? 8'h72 : _GEN_1053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1055 = 8'h1f == io_data_in[47:40] ? 8'hc0 : _GEN_1054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1056 = 8'h20 == io_data_in[47:40] ? 8'hb7 : _GEN_1055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1057 = 8'h21 == io_data_in[47:40] ? 8'hfd : _GEN_1056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1058 = 8'h22 == io_data_in[47:40] ? 8'h93 : _GEN_1057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1059 = 8'h23 == io_data_in[47:40] ? 8'h26 : _GEN_1058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1060 = 8'h24 == io_data_in[47:40] ? 8'h36 : _GEN_1059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1061 = 8'h25 == io_data_in[47:40] ? 8'h3f : _GEN_1060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1062 = 8'h26 == io_data_in[47:40] ? 8'hf7 : _GEN_1061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1063 = 8'h27 == io_data_in[47:40] ? 8'hcc : _GEN_1062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1064 = 8'h28 == io_data_in[47:40] ? 8'h34 : _GEN_1063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1065 = 8'h29 == io_data_in[47:40] ? 8'ha5 : _GEN_1064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1066 = 8'h2a == io_data_in[47:40] ? 8'he5 : _GEN_1065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1067 = 8'h2b == io_data_in[47:40] ? 8'hf1 : _GEN_1066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1068 = 8'h2c == io_data_in[47:40] ? 8'h71 : _GEN_1067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1069 = 8'h2d == io_data_in[47:40] ? 8'hd8 : _GEN_1068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1070 = 8'h2e == io_data_in[47:40] ? 8'h31 : _GEN_1069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1071 = 8'h2f == io_data_in[47:40] ? 8'h15 : _GEN_1070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1072 = 8'h30 == io_data_in[47:40] ? 8'h4 : _GEN_1071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1073 = 8'h31 == io_data_in[47:40] ? 8'hc7 : _GEN_1072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1074 = 8'h32 == io_data_in[47:40] ? 8'h23 : _GEN_1073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1075 = 8'h33 == io_data_in[47:40] ? 8'hc3 : _GEN_1074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1076 = 8'h34 == io_data_in[47:40] ? 8'h18 : _GEN_1075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1077 = 8'h35 == io_data_in[47:40] ? 8'h96 : _GEN_1076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1078 = 8'h36 == io_data_in[47:40] ? 8'h5 : _GEN_1077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1079 = 8'h37 == io_data_in[47:40] ? 8'h9a : _GEN_1078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1080 = 8'h38 == io_data_in[47:40] ? 8'h7 : _GEN_1079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1081 = 8'h39 == io_data_in[47:40] ? 8'h12 : _GEN_1080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1082 = 8'h3a == io_data_in[47:40] ? 8'h80 : _GEN_1081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1083 = 8'h3b == io_data_in[47:40] ? 8'he2 : _GEN_1082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1084 = 8'h3c == io_data_in[47:40] ? 8'heb : _GEN_1083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1085 = 8'h3d == io_data_in[47:40] ? 8'h27 : _GEN_1084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1086 = 8'h3e == io_data_in[47:40] ? 8'hb2 : _GEN_1085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1087 = 8'h3f == io_data_in[47:40] ? 8'h75 : _GEN_1086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1088 = 8'h40 == io_data_in[47:40] ? 8'h9 : _GEN_1087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1089 = 8'h41 == io_data_in[47:40] ? 8'h83 : _GEN_1088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1090 = 8'h42 == io_data_in[47:40] ? 8'h2c : _GEN_1089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1091 = 8'h43 == io_data_in[47:40] ? 8'h1a : _GEN_1090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1092 = 8'h44 == io_data_in[47:40] ? 8'h1b : _GEN_1091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1093 = 8'h45 == io_data_in[47:40] ? 8'h6e : _GEN_1092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1094 = 8'h46 == io_data_in[47:40] ? 8'h5a : _GEN_1093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1095 = 8'h47 == io_data_in[47:40] ? 8'ha0 : _GEN_1094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1096 = 8'h48 == io_data_in[47:40] ? 8'h52 : _GEN_1095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1097 = 8'h49 == io_data_in[47:40] ? 8'h3b : _GEN_1096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1098 = 8'h4a == io_data_in[47:40] ? 8'hd6 : _GEN_1097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1099 = 8'h4b == io_data_in[47:40] ? 8'hb3 : _GEN_1098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1100 = 8'h4c == io_data_in[47:40] ? 8'h29 : _GEN_1099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1101 = 8'h4d == io_data_in[47:40] ? 8'he3 : _GEN_1100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1102 = 8'h4e == io_data_in[47:40] ? 8'h2f : _GEN_1101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1103 = 8'h4f == io_data_in[47:40] ? 8'h84 : _GEN_1102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1104 = 8'h50 == io_data_in[47:40] ? 8'h53 : _GEN_1103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1105 = 8'h51 == io_data_in[47:40] ? 8'hd1 : _GEN_1104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1106 = 8'h52 == io_data_in[47:40] ? 8'h0 : _GEN_1105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1107 = 8'h53 == io_data_in[47:40] ? 8'hed : _GEN_1106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1108 = 8'h54 == io_data_in[47:40] ? 8'h20 : _GEN_1107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1109 = 8'h55 == io_data_in[47:40] ? 8'hfc : _GEN_1108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1110 = 8'h56 == io_data_in[47:40] ? 8'hb1 : _GEN_1109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1111 = 8'h57 == io_data_in[47:40] ? 8'h5b : _GEN_1110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1112 = 8'h58 == io_data_in[47:40] ? 8'h6a : _GEN_1111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1113 = 8'h59 == io_data_in[47:40] ? 8'hcb : _GEN_1112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1114 = 8'h5a == io_data_in[47:40] ? 8'hbe : _GEN_1113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1115 = 8'h5b == io_data_in[47:40] ? 8'h39 : _GEN_1114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1116 = 8'h5c == io_data_in[47:40] ? 8'h4a : _GEN_1115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1117 = 8'h5d == io_data_in[47:40] ? 8'h4c : _GEN_1116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1118 = 8'h5e == io_data_in[47:40] ? 8'h58 : _GEN_1117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1119 = 8'h5f == io_data_in[47:40] ? 8'hcf : _GEN_1118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1120 = 8'h60 == io_data_in[47:40] ? 8'hd0 : _GEN_1119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1121 = 8'h61 == io_data_in[47:40] ? 8'hef : _GEN_1120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1122 = 8'h62 == io_data_in[47:40] ? 8'haa : _GEN_1121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1123 = 8'h63 == io_data_in[47:40] ? 8'hfb : _GEN_1122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1124 = 8'h64 == io_data_in[47:40] ? 8'h43 : _GEN_1123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1125 = 8'h65 == io_data_in[47:40] ? 8'h4d : _GEN_1124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1126 = 8'h66 == io_data_in[47:40] ? 8'h33 : _GEN_1125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1127 = 8'h67 == io_data_in[47:40] ? 8'h85 : _GEN_1126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1128 = 8'h68 == io_data_in[47:40] ? 8'h45 : _GEN_1127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1129 = 8'h69 == io_data_in[47:40] ? 8'hf9 : _GEN_1128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1130 = 8'h6a == io_data_in[47:40] ? 8'h2 : _GEN_1129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1131 = 8'h6b == io_data_in[47:40] ? 8'h7f : _GEN_1130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1132 = 8'h6c == io_data_in[47:40] ? 8'h50 : _GEN_1131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1133 = 8'h6d == io_data_in[47:40] ? 8'h3c : _GEN_1132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1134 = 8'h6e == io_data_in[47:40] ? 8'h9f : _GEN_1133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1135 = 8'h6f == io_data_in[47:40] ? 8'ha8 : _GEN_1134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1136 = 8'h70 == io_data_in[47:40] ? 8'h51 : _GEN_1135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1137 = 8'h71 == io_data_in[47:40] ? 8'ha3 : _GEN_1136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1138 = 8'h72 == io_data_in[47:40] ? 8'h40 : _GEN_1137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1139 = 8'h73 == io_data_in[47:40] ? 8'h8f : _GEN_1138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1140 = 8'h74 == io_data_in[47:40] ? 8'h92 : _GEN_1139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1141 = 8'h75 == io_data_in[47:40] ? 8'h9d : _GEN_1140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1142 = 8'h76 == io_data_in[47:40] ? 8'h38 : _GEN_1141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1143 = 8'h77 == io_data_in[47:40] ? 8'hf5 : _GEN_1142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1144 = 8'h78 == io_data_in[47:40] ? 8'hbc : _GEN_1143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1145 = 8'h79 == io_data_in[47:40] ? 8'hb6 : _GEN_1144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1146 = 8'h7a == io_data_in[47:40] ? 8'hda : _GEN_1145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1147 = 8'h7b == io_data_in[47:40] ? 8'h21 : _GEN_1146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1148 = 8'h7c == io_data_in[47:40] ? 8'h10 : _GEN_1147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1149 = 8'h7d == io_data_in[47:40] ? 8'hff : _GEN_1148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1150 = 8'h7e == io_data_in[47:40] ? 8'hf3 : _GEN_1149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1151 = 8'h7f == io_data_in[47:40] ? 8'hd2 : _GEN_1150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1152 = 8'h80 == io_data_in[47:40] ? 8'hcd : _GEN_1151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1153 = 8'h81 == io_data_in[47:40] ? 8'hc : _GEN_1152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1154 = 8'h82 == io_data_in[47:40] ? 8'h13 : _GEN_1153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1155 = 8'h83 == io_data_in[47:40] ? 8'hec : _GEN_1154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1156 = 8'h84 == io_data_in[47:40] ? 8'h5f : _GEN_1155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1157 = 8'h85 == io_data_in[47:40] ? 8'h97 : _GEN_1156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1158 = 8'h86 == io_data_in[47:40] ? 8'h44 : _GEN_1157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1159 = 8'h87 == io_data_in[47:40] ? 8'h17 : _GEN_1158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1160 = 8'h88 == io_data_in[47:40] ? 8'hc4 : _GEN_1159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1161 = 8'h89 == io_data_in[47:40] ? 8'ha7 : _GEN_1160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1162 = 8'h8a == io_data_in[47:40] ? 8'h7e : _GEN_1161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1163 = 8'h8b == io_data_in[47:40] ? 8'h3d : _GEN_1162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1164 = 8'h8c == io_data_in[47:40] ? 8'h64 : _GEN_1163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1165 = 8'h8d == io_data_in[47:40] ? 8'h5d : _GEN_1164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1166 = 8'h8e == io_data_in[47:40] ? 8'h19 : _GEN_1165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1167 = 8'h8f == io_data_in[47:40] ? 8'h73 : _GEN_1166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1168 = 8'h90 == io_data_in[47:40] ? 8'h60 : _GEN_1167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1169 = 8'h91 == io_data_in[47:40] ? 8'h81 : _GEN_1168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1170 = 8'h92 == io_data_in[47:40] ? 8'h4f : _GEN_1169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1171 = 8'h93 == io_data_in[47:40] ? 8'hdc : _GEN_1170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1172 = 8'h94 == io_data_in[47:40] ? 8'h22 : _GEN_1171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1173 = 8'h95 == io_data_in[47:40] ? 8'h2a : _GEN_1172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1174 = 8'h96 == io_data_in[47:40] ? 8'h90 : _GEN_1173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1175 = 8'h97 == io_data_in[47:40] ? 8'h88 : _GEN_1174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1176 = 8'h98 == io_data_in[47:40] ? 8'h46 : _GEN_1175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1177 = 8'h99 == io_data_in[47:40] ? 8'hee : _GEN_1176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1178 = 8'h9a == io_data_in[47:40] ? 8'hb8 : _GEN_1177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1179 = 8'h9b == io_data_in[47:40] ? 8'h14 : _GEN_1178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1180 = 8'h9c == io_data_in[47:40] ? 8'hde : _GEN_1179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1181 = 8'h9d == io_data_in[47:40] ? 8'h5e : _GEN_1180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1182 = 8'h9e == io_data_in[47:40] ? 8'hb : _GEN_1181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1183 = 8'h9f == io_data_in[47:40] ? 8'hdb : _GEN_1182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1184 = 8'ha0 == io_data_in[47:40] ? 8'he0 : _GEN_1183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1185 = 8'ha1 == io_data_in[47:40] ? 8'h32 : _GEN_1184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1186 = 8'ha2 == io_data_in[47:40] ? 8'h3a : _GEN_1185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1187 = 8'ha3 == io_data_in[47:40] ? 8'ha : _GEN_1186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1188 = 8'ha4 == io_data_in[47:40] ? 8'h49 : _GEN_1187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1189 = 8'ha5 == io_data_in[47:40] ? 8'h6 : _GEN_1188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1190 = 8'ha6 == io_data_in[47:40] ? 8'h24 : _GEN_1189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1191 = 8'ha7 == io_data_in[47:40] ? 8'h5c : _GEN_1190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1192 = 8'ha8 == io_data_in[47:40] ? 8'hc2 : _GEN_1191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1193 = 8'ha9 == io_data_in[47:40] ? 8'hd3 : _GEN_1192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1194 = 8'haa == io_data_in[47:40] ? 8'hac : _GEN_1193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1195 = 8'hab == io_data_in[47:40] ? 8'h62 : _GEN_1194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1196 = 8'hac == io_data_in[47:40] ? 8'h91 : _GEN_1195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1197 = 8'had == io_data_in[47:40] ? 8'h95 : _GEN_1196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1198 = 8'hae == io_data_in[47:40] ? 8'he4 : _GEN_1197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1199 = 8'haf == io_data_in[47:40] ? 8'h79 : _GEN_1198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1200 = 8'hb0 == io_data_in[47:40] ? 8'he7 : _GEN_1199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1201 = 8'hb1 == io_data_in[47:40] ? 8'hc8 : _GEN_1200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1202 = 8'hb2 == io_data_in[47:40] ? 8'h37 : _GEN_1201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1203 = 8'hb3 == io_data_in[47:40] ? 8'h6d : _GEN_1202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1204 = 8'hb4 == io_data_in[47:40] ? 8'h8d : _GEN_1203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1205 = 8'hb5 == io_data_in[47:40] ? 8'hd5 : _GEN_1204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1206 = 8'hb6 == io_data_in[47:40] ? 8'h4e : _GEN_1205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1207 = 8'hb7 == io_data_in[47:40] ? 8'ha9 : _GEN_1206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1208 = 8'hb8 == io_data_in[47:40] ? 8'h6c : _GEN_1207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1209 = 8'hb9 == io_data_in[47:40] ? 8'h56 : _GEN_1208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1210 = 8'hba == io_data_in[47:40] ? 8'hf4 : _GEN_1209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1211 = 8'hbb == io_data_in[47:40] ? 8'hea : _GEN_1210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1212 = 8'hbc == io_data_in[47:40] ? 8'h65 : _GEN_1211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1213 = 8'hbd == io_data_in[47:40] ? 8'h7a : _GEN_1212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1214 = 8'hbe == io_data_in[47:40] ? 8'hae : _GEN_1213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1215 = 8'hbf == io_data_in[47:40] ? 8'h8 : _GEN_1214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1216 = 8'hc0 == io_data_in[47:40] ? 8'hba : _GEN_1215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1217 = 8'hc1 == io_data_in[47:40] ? 8'h78 : _GEN_1216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1218 = 8'hc2 == io_data_in[47:40] ? 8'h25 : _GEN_1217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1219 = 8'hc3 == io_data_in[47:40] ? 8'h2e : _GEN_1218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1220 = 8'hc4 == io_data_in[47:40] ? 8'h1c : _GEN_1219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1221 = 8'hc5 == io_data_in[47:40] ? 8'ha6 : _GEN_1220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1222 = 8'hc6 == io_data_in[47:40] ? 8'hb4 : _GEN_1221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1223 = 8'hc7 == io_data_in[47:40] ? 8'hc6 : _GEN_1222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1224 = 8'hc8 == io_data_in[47:40] ? 8'he8 : _GEN_1223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1225 = 8'hc9 == io_data_in[47:40] ? 8'hdd : _GEN_1224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1226 = 8'hca == io_data_in[47:40] ? 8'h74 : _GEN_1225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1227 = 8'hcb == io_data_in[47:40] ? 8'h1f : _GEN_1226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1228 = 8'hcc == io_data_in[47:40] ? 8'h4b : _GEN_1227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1229 = 8'hcd == io_data_in[47:40] ? 8'hbd : _GEN_1228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1230 = 8'hce == io_data_in[47:40] ? 8'h8b : _GEN_1229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1231 = 8'hcf == io_data_in[47:40] ? 8'h8a : _GEN_1230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1232 = 8'hd0 == io_data_in[47:40] ? 8'h70 : _GEN_1231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1233 = 8'hd1 == io_data_in[47:40] ? 8'h3e : _GEN_1232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1234 = 8'hd2 == io_data_in[47:40] ? 8'hb5 : _GEN_1233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1235 = 8'hd3 == io_data_in[47:40] ? 8'h66 : _GEN_1234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1236 = 8'hd4 == io_data_in[47:40] ? 8'h48 : _GEN_1235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1237 = 8'hd5 == io_data_in[47:40] ? 8'h3 : _GEN_1236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1238 = 8'hd6 == io_data_in[47:40] ? 8'hf6 : _GEN_1237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1239 = 8'hd7 == io_data_in[47:40] ? 8'he : _GEN_1238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1240 = 8'hd8 == io_data_in[47:40] ? 8'h61 : _GEN_1239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1241 = 8'hd9 == io_data_in[47:40] ? 8'h35 : _GEN_1240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1242 = 8'hda == io_data_in[47:40] ? 8'h57 : _GEN_1241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1243 = 8'hdb == io_data_in[47:40] ? 8'hb9 : _GEN_1242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1244 = 8'hdc == io_data_in[47:40] ? 8'h86 : _GEN_1243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1245 = 8'hdd == io_data_in[47:40] ? 8'hc1 : _GEN_1244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1246 = 8'hde == io_data_in[47:40] ? 8'h1d : _GEN_1245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1247 = 8'hdf == io_data_in[47:40] ? 8'h9e : _GEN_1246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1248 = 8'he0 == io_data_in[47:40] ? 8'he1 : _GEN_1247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1249 = 8'he1 == io_data_in[47:40] ? 8'hf8 : _GEN_1248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1250 = 8'he2 == io_data_in[47:40] ? 8'h98 : _GEN_1249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1251 = 8'he3 == io_data_in[47:40] ? 8'h11 : _GEN_1250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1252 = 8'he4 == io_data_in[47:40] ? 8'h69 : _GEN_1251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1253 = 8'he5 == io_data_in[47:40] ? 8'hd9 : _GEN_1252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1254 = 8'he6 == io_data_in[47:40] ? 8'h8e : _GEN_1253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1255 = 8'he7 == io_data_in[47:40] ? 8'h94 : _GEN_1254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1256 = 8'he8 == io_data_in[47:40] ? 8'h9b : _GEN_1255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1257 = 8'he9 == io_data_in[47:40] ? 8'h1e : _GEN_1256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1258 = 8'hea == io_data_in[47:40] ? 8'h87 : _GEN_1257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1259 = 8'heb == io_data_in[47:40] ? 8'he9 : _GEN_1258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1260 = 8'hec == io_data_in[47:40] ? 8'hce : _GEN_1259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1261 = 8'hed == io_data_in[47:40] ? 8'h55 : _GEN_1260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1262 = 8'hee == io_data_in[47:40] ? 8'h28 : _GEN_1261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1263 = 8'hef == io_data_in[47:40] ? 8'hdf : _GEN_1262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1264 = 8'hf0 == io_data_in[47:40] ? 8'h8c : _GEN_1263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1265 = 8'hf1 == io_data_in[47:40] ? 8'ha1 : _GEN_1264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1266 = 8'hf2 == io_data_in[47:40] ? 8'h89 : _GEN_1265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1267 = 8'hf3 == io_data_in[47:40] ? 8'hd : _GEN_1266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1268 = 8'hf4 == io_data_in[47:40] ? 8'hbf : _GEN_1267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1269 = 8'hf5 == io_data_in[47:40] ? 8'he6 : _GEN_1268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1270 = 8'hf6 == io_data_in[47:40] ? 8'h42 : _GEN_1269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1271 = 8'hf7 == io_data_in[47:40] ? 8'h68 : _GEN_1270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1272 = 8'hf8 == io_data_in[47:40] ? 8'h41 : _GEN_1271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1273 = 8'hf9 == io_data_in[47:40] ? 8'h99 : _GEN_1272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1274 = 8'hfa == io_data_in[47:40] ? 8'h2d : _GEN_1273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1275 = 8'hfb == io_data_in[47:40] ? 8'hf : _GEN_1274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1276 = 8'hfc == io_data_in[47:40] ? 8'hb0 : _GEN_1275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1277 = 8'hfd == io_data_in[47:40] ? 8'h54 : _GEN_1276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1278 = 8'hfe == io_data_in[47:40] ? 8'hbb : _GEN_1277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1279 = 8'hff == io_data_in[47:40] ? 8'h16 : _GEN_1278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1281 = 8'h1 == io_data_in[39:32] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1282 = 8'h2 == io_data_in[39:32] ? 8'h77 : _GEN_1281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1283 = 8'h3 == io_data_in[39:32] ? 8'h7b : _GEN_1282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1284 = 8'h4 == io_data_in[39:32] ? 8'hf2 : _GEN_1283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1285 = 8'h5 == io_data_in[39:32] ? 8'h6b : _GEN_1284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1286 = 8'h6 == io_data_in[39:32] ? 8'h6f : _GEN_1285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1287 = 8'h7 == io_data_in[39:32] ? 8'hc5 : _GEN_1286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1288 = 8'h8 == io_data_in[39:32] ? 8'h30 : _GEN_1287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1289 = 8'h9 == io_data_in[39:32] ? 8'h1 : _GEN_1288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1290 = 8'ha == io_data_in[39:32] ? 8'h67 : _GEN_1289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1291 = 8'hb == io_data_in[39:32] ? 8'h2b : _GEN_1290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1292 = 8'hc == io_data_in[39:32] ? 8'hfe : _GEN_1291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1293 = 8'hd == io_data_in[39:32] ? 8'hd7 : _GEN_1292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1294 = 8'he == io_data_in[39:32] ? 8'hab : _GEN_1293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1295 = 8'hf == io_data_in[39:32] ? 8'h76 : _GEN_1294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1296 = 8'h10 == io_data_in[39:32] ? 8'hca : _GEN_1295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1297 = 8'h11 == io_data_in[39:32] ? 8'h82 : _GEN_1296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1298 = 8'h12 == io_data_in[39:32] ? 8'hc9 : _GEN_1297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1299 = 8'h13 == io_data_in[39:32] ? 8'h7d : _GEN_1298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1300 = 8'h14 == io_data_in[39:32] ? 8'hfa : _GEN_1299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1301 = 8'h15 == io_data_in[39:32] ? 8'h59 : _GEN_1300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1302 = 8'h16 == io_data_in[39:32] ? 8'h47 : _GEN_1301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1303 = 8'h17 == io_data_in[39:32] ? 8'hf0 : _GEN_1302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1304 = 8'h18 == io_data_in[39:32] ? 8'had : _GEN_1303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1305 = 8'h19 == io_data_in[39:32] ? 8'hd4 : _GEN_1304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1306 = 8'h1a == io_data_in[39:32] ? 8'ha2 : _GEN_1305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1307 = 8'h1b == io_data_in[39:32] ? 8'haf : _GEN_1306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1308 = 8'h1c == io_data_in[39:32] ? 8'h9c : _GEN_1307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1309 = 8'h1d == io_data_in[39:32] ? 8'ha4 : _GEN_1308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1310 = 8'h1e == io_data_in[39:32] ? 8'h72 : _GEN_1309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1311 = 8'h1f == io_data_in[39:32] ? 8'hc0 : _GEN_1310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1312 = 8'h20 == io_data_in[39:32] ? 8'hb7 : _GEN_1311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1313 = 8'h21 == io_data_in[39:32] ? 8'hfd : _GEN_1312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1314 = 8'h22 == io_data_in[39:32] ? 8'h93 : _GEN_1313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1315 = 8'h23 == io_data_in[39:32] ? 8'h26 : _GEN_1314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1316 = 8'h24 == io_data_in[39:32] ? 8'h36 : _GEN_1315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1317 = 8'h25 == io_data_in[39:32] ? 8'h3f : _GEN_1316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1318 = 8'h26 == io_data_in[39:32] ? 8'hf7 : _GEN_1317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1319 = 8'h27 == io_data_in[39:32] ? 8'hcc : _GEN_1318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1320 = 8'h28 == io_data_in[39:32] ? 8'h34 : _GEN_1319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1321 = 8'h29 == io_data_in[39:32] ? 8'ha5 : _GEN_1320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1322 = 8'h2a == io_data_in[39:32] ? 8'he5 : _GEN_1321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1323 = 8'h2b == io_data_in[39:32] ? 8'hf1 : _GEN_1322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1324 = 8'h2c == io_data_in[39:32] ? 8'h71 : _GEN_1323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1325 = 8'h2d == io_data_in[39:32] ? 8'hd8 : _GEN_1324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1326 = 8'h2e == io_data_in[39:32] ? 8'h31 : _GEN_1325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1327 = 8'h2f == io_data_in[39:32] ? 8'h15 : _GEN_1326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1328 = 8'h30 == io_data_in[39:32] ? 8'h4 : _GEN_1327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1329 = 8'h31 == io_data_in[39:32] ? 8'hc7 : _GEN_1328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1330 = 8'h32 == io_data_in[39:32] ? 8'h23 : _GEN_1329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1331 = 8'h33 == io_data_in[39:32] ? 8'hc3 : _GEN_1330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1332 = 8'h34 == io_data_in[39:32] ? 8'h18 : _GEN_1331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1333 = 8'h35 == io_data_in[39:32] ? 8'h96 : _GEN_1332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1334 = 8'h36 == io_data_in[39:32] ? 8'h5 : _GEN_1333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1335 = 8'h37 == io_data_in[39:32] ? 8'h9a : _GEN_1334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1336 = 8'h38 == io_data_in[39:32] ? 8'h7 : _GEN_1335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1337 = 8'h39 == io_data_in[39:32] ? 8'h12 : _GEN_1336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1338 = 8'h3a == io_data_in[39:32] ? 8'h80 : _GEN_1337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1339 = 8'h3b == io_data_in[39:32] ? 8'he2 : _GEN_1338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1340 = 8'h3c == io_data_in[39:32] ? 8'heb : _GEN_1339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1341 = 8'h3d == io_data_in[39:32] ? 8'h27 : _GEN_1340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1342 = 8'h3e == io_data_in[39:32] ? 8'hb2 : _GEN_1341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1343 = 8'h3f == io_data_in[39:32] ? 8'h75 : _GEN_1342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1344 = 8'h40 == io_data_in[39:32] ? 8'h9 : _GEN_1343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1345 = 8'h41 == io_data_in[39:32] ? 8'h83 : _GEN_1344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1346 = 8'h42 == io_data_in[39:32] ? 8'h2c : _GEN_1345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1347 = 8'h43 == io_data_in[39:32] ? 8'h1a : _GEN_1346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1348 = 8'h44 == io_data_in[39:32] ? 8'h1b : _GEN_1347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1349 = 8'h45 == io_data_in[39:32] ? 8'h6e : _GEN_1348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1350 = 8'h46 == io_data_in[39:32] ? 8'h5a : _GEN_1349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1351 = 8'h47 == io_data_in[39:32] ? 8'ha0 : _GEN_1350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1352 = 8'h48 == io_data_in[39:32] ? 8'h52 : _GEN_1351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1353 = 8'h49 == io_data_in[39:32] ? 8'h3b : _GEN_1352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1354 = 8'h4a == io_data_in[39:32] ? 8'hd6 : _GEN_1353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1355 = 8'h4b == io_data_in[39:32] ? 8'hb3 : _GEN_1354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1356 = 8'h4c == io_data_in[39:32] ? 8'h29 : _GEN_1355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1357 = 8'h4d == io_data_in[39:32] ? 8'he3 : _GEN_1356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1358 = 8'h4e == io_data_in[39:32] ? 8'h2f : _GEN_1357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1359 = 8'h4f == io_data_in[39:32] ? 8'h84 : _GEN_1358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1360 = 8'h50 == io_data_in[39:32] ? 8'h53 : _GEN_1359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1361 = 8'h51 == io_data_in[39:32] ? 8'hd1 : _GEN_1360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1362 = 8'h52 == io_data_in[39:32] ? 8'h0 : _GEN_1361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1363 = 8'h53 == io_data_in[39:32] ? 8'hed : _GEN_1362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1364 = 8'h54 == io_data_in[39:32] ? 8'h20 : _GEN_1363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1365 = 8'h55 == io_data_in[39:32] ? 8'hfc : _GEN_1364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1366 = 8'h56 == io_data_in[39:32] ? 8'hb1 : _GEN_1365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1367 = 8'h57 == io_data_in[39:32] ? 8'h5b : _GEN_1366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1368 = 8'h58 == io_data_in[39:32] ? 8'h6a : _GEN_1367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1369 = 8'h59 == io_data_in[39:32] ? 8'hcb : _GEN_1368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1370 = 8'h5a == io_data_in[39:32] ? 8'hbe : _GEN_1369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1371 = 8'h5b == io_data_in[39:32] ? 8'h39 : _GEN_1370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1372 = 8'h5c == io_data_in[39:32] ? 8'h4a : _GEN_1371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1373 = 8'h5d == io_data_in[39:32] ? 8'h4c : _GEN_1372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1374 = 8'h5e == io_data_in[39:32] ? 8'h58 : _GEN_1373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1375 = 8'h5f == io_data_in[39:32] ? 8'hcf : _GEN_1374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1376 = 8'h60 == io_data_in[39:32] ? 8'hd0 : _GEN_1375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1377 = 8'h61 == io_data_in[39:32] ? 8'hef : _GEN_1376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1378 = 8'h62 == io_data_in[39:32] ? 8'haa : _GEN_1377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1379 = 8'h63 == io_data_in[39:32] ? 8'hfb : _GEN_1378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1380 = 8'h64 == io_data_in[39:32] ? 8'h43 : _GEN_1379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1381 = 8'h65 == io_data_in[39:32] ? 8'h4d : _GEN_1380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1382 = 8'h66 == io_data_in[39:32] ? 8'h33 : _GEN_1381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1383 = 8'h67 == io_data_in[39:32] ? 8'h85 : _GEN_1382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1384 = 8'h68 == io_data_in[39:32] ? 8'h45 : _GEN_1383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1385 = 8'h69 == io_data_in[39:32] ? 8'hf9 : _GEN_1384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1386 = 8'h6a == io_data_in[39:32] ? 8'h2 : _GEN_1385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1387 = 8'h6b == io_data_in[39:32] ? 8'h7f : _GEN_1386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1388 = 8'h6c == io_data_in[39:32] ? 8'h50 : _GEN_1387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1389 = 8'h6d == io_data_in[39:32] ? 8'h3c : _GEN_1388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1390 = 8'h6e == io_data_in[39:32] ? 8'h9f : _GEN_1389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1391 = 8'h6f == io_data_in[39:32] ? 8'ha8 : _GEN_1390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1392 = 8'h70 == io_data_in[39:32] ? 8'h51 : _GEN_1391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1393 = 8'h71 == io_data_in[39:32] ? 8'ha3 : _GEN_1392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1394 = 8'h72 == io_data_in[39:32] ? 8'h40 : _GEN_1393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1395 = 8'h73 == io_data_in[39:32] ? 8'h8f : _GEN_1394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1396 = 8'h74 == io_data_in[39:32] ? 8'h92 : _GEN_1395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1397 = 8'h75 == io_data_in[39:32] ? 8'h9d : _GEN_1396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1398 = 8'h76 == io_data_in[39:32] ? 8'h38 : _GEN_1397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1399 = 8'h77 == io_data_in[39:32] ? 8'hf5 : _GEN_1398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1400 = 8'h78 == io_data_in[39:32] ? 8'hbc : _GEN_1399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1401 = 8'h79 == io_data_in[39:32] ? 8'hb6 : _GEN_1400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1402 = 8'h7a == io_data_in[39:32] ? 8'hda : _GEN_1401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1403 = 8'h7b == io_data_in[39:32] ? 8'h21 : _GEN_1402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1404 = 8'h7c == io_data_in[39:32] ? 8'h10 : _GEN_1403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1405 = 8'h7d == io_data_in[39:32] ? 8'hff : _GEN_1404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1406 = 8'h7e == io_data_in[39:32] ? 8'hf3 : _GEN_1405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1407 = 8'h7f == io_data_in[39:32] ? 8'hd2 : _GEN_1406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1408 = 8'h80 == io_data_in[39:32] ? 8'hcd : _GEN_1407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1409 = 8'h81 == io_data_in[39:32] ? 8'hc : _GEN_1408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1410 = 8'h82 == io_data_in[39:32] ? 8'h13 : _GEN_1409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1411 = 8'h83 == io_data_in[39:32] ? 8'hec : _GEN_1410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1412 = 8'h84 == io_data_in[39:32] ? 8'h5f : _GEN_1411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1413 = 8'h85 == io_data_in[39:32] ? 8'h97 : _GEN_1412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1414 = 8'h86 == io_data_in[39:32] ? 8'h44 : _GEN_1413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1415 = 8'h87 == io_data_in[39:32] ? 8'h17 : _GEN_1414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1416 = 8'h88 == io_data_in[39:32] ? 8'hc4 : _GEN_1415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1417 = 8'h89 == io_data_in[39:32] ? 8'ha7 : _GEN_1416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1418 = 8'h8a == io_data_in[39:32] ? 8'h7e : _GEN_1417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1419 = 8'h8b == io_data_in[39:32] ? 8'h3d : _GEN_1418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1420 = 8'h8c == io_data_in[39:32] ? 8'h64 : _GEN_1419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1421 = 8'h8d == io_data_in[39:32] ? 8'h5d : _GEN_1420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1422 = 8'h8e == io_data_in[39:32] ? 8'h19 : _GEN_1421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1423 = 8'h8f == io_data_in[39:32] ? 8'h73 : _GEN_1422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1424 = 8'h90 == io_data_in[39:32] ? 8'h60 : _GEN_1423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1425 = 8'h91 == io_data_in[39:32] ? 8'h81 : _GEN_1424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1426 = 8'h92 == io_data_in[39:32] ? 8'h4f : _GEN_1425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1427 = 8'h93 == io_data_in[39:32] ? 8'hdc : _GEN_1426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1428 = 8'h94 == io_data_in[39:32] ? 8'h22 : _GEN_1427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1429 = 8'h95 == io_data_in[39:32] ? 8'h2a : _GEN_1428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1430 = 8'h96 == io_data_in[39:32] ? 8'h90 : _GEN_1429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1431 = 8'h97 == io_data_in[39:32] ? 8'h88 : _GEN_1430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1432 = 8'h98 == io_data_in[39:32] ? 8'h46 : _GEN_1431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1433 = 8'h99 == io_data_in[39:32] ? 8'hee : _GEN_1432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1434 = 8'h9a == io_data_in[39:32] ? 8'hb8 : _GEN_1433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1435 = 8'h9b == io_data_in[39:32] ? 8'h14 : _GEN_1434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1436 = 8'h9c == io_data_in[39:32] ? 8'hde : _GEN_1435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1437 = 8'h9d == io_data_in[39:32] ? 8'h5e : _GEN_1436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1438 = 8'h9e == io_data_in[39:32] ? 8'hb : _GEN_1437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1439 = 8'h9f == io_data_in[39:32] ? 8'hdb : _GEN_1438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1440 = 8'ha0 == io_data_in[39:32] ? 8'he0 : _GEN_1439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1441 = 8'ha1 == io_data_in[39:32] ? 8'h32 : _GEN_1440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1442 = 8'ha2 == io_data_in[39:32] ? 8'h3a : _GEN_1441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1443 = 8'ha3 == io_data_in[39:32] ? 8'ha : _GEN_1442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1444 = 8'ha4 == io_data_in[39:32] ? 8'h49 : _GEN_1443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1445 = 8'ha5 == io_data_in[39:32] ? 8'h6 : _GEN_1444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1446 = 8'ha6 == io_data_in[39:32] ? 8'h24 : _GEN_1445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1447 = 8'ha7 == io_data_in[39:32] ? 8'h5c : _GEN_1446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1448 = 8'ha8 == io_data_in[39:32] ? 8'hc2 : _GEN_1447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1449 = 8'ha9 == io_data_in[39:32] ? 8'hd3 : _GEN_1448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1450 = 8'haa == io_data_in[39:32] ? 8'hac : _GEN_1449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1451 = 8'hab == io_data_in[39:32] ? 8'h62 : _GEN_1450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1452 = 8'hac == io_data_in[39:32] ? 8'h91 : _GEN_1451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1453 = 8'had == io_data_in[39:32] ? 8'h95 : _GEN_1452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1454 = 8'hae == io_data_in[39:32] ? 8'he4 : _GEN_1453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1455 = 8'haf == io_data_in[39:32] ? 8'h79 : _GEN_1454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1456 = 8'hb0 == io_data_in[39:32] ? 8'he7 : _GEN_1455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1457 = 8'hb1 == io_data_in[39:32] ? 8'hc8 : _GEN_1456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1458 = 8'hb2 == io_data_in[39:32] ? 8'h37 : _GEN_1457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1459 = 8'hb3 == io_data_in[39:32] ? 8'h6d : _GEN_1458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1460 = 8'hb4 == io_data_in[39:32] ? 8'h8d : _GEN_1459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1461 = 8'hb5 == io_data_in[39:32] ? 8'hd5 : _GEN_1460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1462 = 8'hb6 == io_data_in[39:32] ? 8'h4e : _GEN_1461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1463 = 8'hb7 == io_data_in[39:32] ? 8'ha9 : _GEN_1462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1464 = 8'hb8 == io_data_in[39:32] ? 8'h6c : _GEN_1463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1465 = 8'hb9 == io_data_in[39:32] ? 8'h56 : _GEN_1464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1466 = 8'hba == io_data_in[39:32] ? 8'hf4 : _GEN_1465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1467 = 8'hbb == io_data_in[39:32] ? 8'hea : _GEN_1466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1468 = 8'hbc == io_data_in[39:32] ? 8'h65 : _GEN_1467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1469 = 8'hbd == io_data_in[39:32] ? 8'h7a : _GEN_1468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1470 = 8'hbe == io_data_in[39:32] ? 8'hae : _GEN_1469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1471 = 8'hbf == io_data_in[39:32] ? 8'h8 : _GEN_1470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1472 = 8'hc0 == io_data_in[39:32] ? 8'hba : _GEN_1471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1473 = 8'hc1 == io_data_in[39:32] ? 8'h78 : _GEN_1472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1474 = 8'hc2 == io_data_in[39:32] ? 8'h25 : _GEN_1473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1475 = 8'hc3 == io_data_in[39:32] ? 8'h2e : _GEN_1474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1476 = 8'hc4 == io_data_in[39:32] ? 8'h1c : _GEN_1475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1477 = 8'hc5 == io_data_in[39:32] ? 8'ha6 : _GEN_1476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1478 = 8'hc6 == io_data_in[39:32] ? 8'hb4 : _GEN_1477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1479 = 8'hc7 == io_data_in[39:32] ? 8'hc6 : _GEN_1478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1480 = 8'hc8 == io_data_in[39:32] ? 8'he8 : _GEN_1479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1481 = 8'hc9 == io_data_in[39:32] ? 8'hdd : _GEN_1480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1482 = 8'hca == io_data_in[39:32] ? 8'h74 : _GEN_1481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1483 = 8'hcb == io_data_in[39:32] ? 8'h1f : _GEN_1482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1484 = 8'hcc == io_data_in[39:32] ? 8'h4b : _GEN_1483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1485 = 8'hcd == io_data_in[39:32] ? 8'hbd : _GEN_1484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1486 = 8'hce == io_data_in[39:32] ? 8'h8b : _GEN_1485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1487 = 8'hcf == io_data_in[39:32] ? 8'h8a : _GEN_1486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1488 = 8'hd0 == io_data_in[39:32] ? 8'h70 : _GEN_1487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1489 = 8'hd1 == io_data_in[39:32] ? 8'h3e : _GEN_1488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1490 = 8'hd2 == io_data_in[39:32] ? 8'hb5 : _GEN_1489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1491 = 8'hd3 == io_data_in[39:32] ? 8'h66 : _GEN_1490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1492 = 8'hd4 == io_data_in[39:32] ? 8'h48 : _GEN_1491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1493 = 8'hd5 == io_data_in[39:32] ? 8'h3 : _GEN_1492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1494 = 8'hd6 == io_data_in[39:32] ? 8'hf6 : _GEN_1493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1495 = 8'hd7 == io_data_in[39:32] ? 8'he : _GEN_1494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1496 = 8'hd8 == io_data_in[39:32] ? 8'h61 : _GEN_1495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1497 = 8'hd9 == io_data_in[39:32] ? 8'h35 : _GEN_1496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1498 = 8'hda == io_data_in[39:32] ? 8'h57 : _GEN_1497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1499 = 8'hdb == io_data_in[39:32] ? 8'hb9 : _GEN_1498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1500 = 8'hdc == io_data_in[39:32] ? 8'h86 : _GEN_1499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1501 = 8'hdd == io_data_in[39:32] ? 8'hc1 : _GEN_1500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1502 = 8'hde == io_data_in[39:32] ? 8'h1d : _GEN_1501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1503 = 8'hdf == io_data_in[39:32] ? 8'h9e : _GEN_1502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1504 = 8'he0 == io_data_in[39:32] ? 8'he1 : _GEN_1503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1505 = 8'he1 == io_data_in[39:32] ? 8'hf8 : _GEN_1504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1506 = 8'he2 == io_data_in[39:32] ? 8'h98 : _GEN_1505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1507 = 8'he3 == io_data_in[39:32] ? 8'h11 : _GEN_1506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1508 = 8'he4 == io_data_in[39:32] ? 8'h69 : _GEN_1507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1509 = 8'he5 == io_data_in[39:32] ? 8'hd9 : _GEN_1508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1510 = 8'he6 == io_data_in[39:32] ? 8'h8e : _GEN_1509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1511 = 8'he7 == io_data_in[39:32] ? 8'h94 : _GEN_1510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1512 = 8'he8 == io_data_in[39:32] ? 8'h9b : _GEN_1511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1513 = 8'he9 == io_data_in[39:32] ? 8'h1e : _GEN_1512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1514 = 8'hea == io_data_in[39:32] ? 8'h87 : _GEN_1513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1515 = 8'heb == io_data_in[39:32] ? 8'he9 : _GEN_1514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1516 = 8'hec == io_data_in[39:32] ? 8'hce : _GEN_1515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1517 = 8'hed == io_data_in[39:32] ? 8'h55 : _GEN_1516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1518 = 8'hee == io_data_in[39:32] ? 8'h28 : _GEN_1517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1519 = 8'hef == io_data_in[39:32] ? 8'hdf : _GEN_1518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1520 = 8'hf0 == io_data_in[39:32] ? 8'h8c : _GEN_1519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1521 = 8'hf1 == io_data_in[39:32] ? 8'ha1 : _GEN_1520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1522 = 8'hf2 == io_data_in[39:32] ? 8'h89 : _GEN_1521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1523 = 8'hf3 == io_data_in[39:32] ? 8'hd : _GEN_1522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1524 = 8'hf4 == io_data_in[39:32] ? 8'hbf : _GEN_1523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1525 = 8'hf5 == io_data_in[39:32] ? 8'he6 : _GEN_1524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1526 = 8'hf6 == io_data_in[39:32] ? 8'h42 : _GEN_1525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1527 = 8'hf7 == io_data_in[39:32] ? 8'h68 : _GEN_1526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1528 = 8'hf8 == io_data_in[39:32] ? 8'h41 : _GEN_1527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1529 = 8'hf9 == io_data_in[39:32] ? 8'h99 : _GEN_1528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1530 = 8'hfa == io_data_in[39:32] ? 8'h2d : _GEN_1529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1531 = 8'hfb == io_data_in[39:32] ? 8'hf : _GEN_1530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1532 = 8'hfc == io_data_in[39:32] ? 8'hb0 : _GEN_1531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1533 = 8'hfd == io_data_in[39:32] ? 8'h54 : _GEN_1532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1534 = 8'hfe == io_data_in[39:32] ? 8'hbb : _GEN_1533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1535 = 8'hff == io_data_in[39:32] ? 8'h16 : _GEN_1534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1537 = 8'h1 == io_data_in[63:56] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1538 = 8'h2 == io_data_in[63:56] ? 8'h77 : _GEN_1537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1539 = 8'h3 == io_data_in[63:56] ? 8'h7b : _GEN_1538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1540 = 8'h4 == io_data_in[63:56] ? 8'hf2 : _GEN_1539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1541 = 8'h5 == io_data_in[63:56] ? 8'h6b : _GEN_1540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1542 = 8'h6 == io_data_in[63:56] ? 8'h6f : _GEN_1541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1543 = 8'h7 == io_data_in[63:56] ? 8'hc5 : _GEN_1542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1544 = 8'h8 == io_data_in[63:56] ? 8'h30 : _GEN_1543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1545 = 8'h9 == io_data_in[63:56] ? 8'h1 : _GEN_1544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1546 = 8'ha == io_data_in[63:56] ? 8'h67 : _GEN_1545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1547 = 8'hb == io_data_in[63:56] ? 8'h2b : _GEN_1546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1548 = 8'hc == io_data_in[63:56] ? 8'hfe : _GEN_1547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1549 = 8'hd == io_data_in[63:56] ? 8'hd7 : _GEN_1548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1550 = 8'he == io_data_in[63:56] ? 8'hab : _GEN_1549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1551 = 8'hf == io_data_in[63:56] ? 8'h76 : _GEN_1550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1552 = 8'h10 == io_data_in[63:56] ? 8'hca : _GEN_1551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1553 = 8'h11 == io_data_in[63:56] ? 8'h82 : _GEN_1552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1554 = 8'h12 == io_data_in[63:56] ? 8'hc9 : _GEN_1553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1555 = 8'h13 == io_data_in[63:56] ? 8'h7d : _GEN_1554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1556 = 8'h14 == io_data_in[63:56] ? 8'hfa : _GEN_1555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1557 = 8'h15 == io_data_in[63:56] ? 8'h59 : _GEN_1556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1558 = 8'h16 == io_data_in[63:56] ? 8'h47 : _GEN_1557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1559 = 8'h17 == io_data_in[63:56] ? 8'hf0 : _GEN_1558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1560 = 8'h18 == io_data_in[63:56] ? 8'had : _GEN_1559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1561 = 8'h19 == io_data_in[63:56] ? 8'hd4 : _GEN_1560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1562 = 8'h1a == io_data_in[63:56] ? 8'ha2 : _GEN_1561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1563 = 8'h1b == io_data_in[63:56] ? 8'haf : _GEN_1562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1564 = 8'h1c == io_data_in[63:56] ? 8'h9c : _GEN_1563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1565 = 8'h1d == io_data_in[63:56] ? 8'ha4 : _GEN_1564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1566 = 8'h1e == io_data_in[63:56] ? 8'h72 : _GEN_1565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1567 = 8'h1f == io_data_in[63:56] ? 8'hc0 : _GEN_1566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1568 = 8'h20 == io_data_in[63:56] ? 8'hb7 : _GEN_1567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1569 = 8'h21 == io_data_in[63:56] ? 8'hfd : _GEN_1568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1570 = 8'h22 == io_data_in[63:56] ? 8'h93 : _GEN_1569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1571 = 8'h23 == io_data_in[63:56] ? 8'h26 : _GEN_1570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1572 = 8'h24 == io_data_in[63:56] ? 8'h36 : _GEN_1571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1573 = 8'h25 == io_data_in[63:56] ? 8'h3f : _GEN_1572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1574 = 8'h26 == io_data_in[63:56] ? 8'hf7 : _GEN_1573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1575 = 8'h27 == io_data_in[63:56] ? 8'hcc : _GEN_1574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1576 = 8'h28 == io_data_in[63:56] ? 8'h34 : _GEN_1575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1577 = 8'h29 == io_data_in[63:56] ? 8'ha5 : _GEN_1576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1578 = 8'h2a == io_data_in[63:56] ? 8'he5 : _GEN_1577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1579 = 8'h2b == io_data_in[63:56] ? 8'hf1 : _GEN_1578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1580 = 8'h2c == io_data_in[63:56] ? 8'h71 : _GEN_1579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1581 = 8'h2d == io_data_in[63:56] ? 8'hd8 : _GEN_1580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1582 = 8'h2e == io_data_in[63:56] ? 8'h31 : _GEN_1581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1583 = 8'h2f == io_data_in[63:56] ? 8'h15 : _GEN_1582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1584 = 8'h30 == io_data_in[63:56] ? 8'h4 : _GEN_1583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1585 = 8'h31 == io_data_in[63:56] ? 8'hc7 : _GEN_1584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1586 = 8'h32 == io_data_in[63:56] ? 8'h23 : _GEN_1585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1587 = 8'h33 == io_data_in[63:56] ? 8'hc3 : _GEN_1586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1588 = 8'h34 == io_data_in[63:56] ? 8'h18 : _GEN_1587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1589 = 8'h35 == io_data_in[63:56] ? 8'h96 : _GEN_1588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1590 = 8'h36 == io_data_in[63:56] ? 8'h5 : _GEN_1589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1591 = 8'h37 == io_data_in[63:56] ? 8'h9a : _GEN_1590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1592 = 8'h38 == io_data_in[63:56] ? 8'h7 : _GEN_1591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1593 = 8'h39 == io_data_in[63:56] ? 8'h12 : _GEN_1592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1594 = 8'h3a == io_data_in[63:56] ? 8'h80 : _GEN_1593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1595 = 8'h3b == io_data_in[63:56] ? 8'he2 : _GEN_1594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1596 = 8'h3c == io_data_in[63:56] ? 8'heb : _GEN_1595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1597 = 8'h3d == io_data_in[63:56] ? 8'h27 : _GEN_1596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1598 = 8'h3e == io_data_in[63:56] ? 8'hb2 : _GEN_1597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1599 = 8'h3f == io_data_in[63:56] ? 8'h75 : _GEN_1598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1600 = 8'h40 == io_data_in[63:56] ? 8'h9 : _GEN_1599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1601 = 8'h41 == io_data_in[63:56] ? 8'h83 : _GEN_1600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1602 = 8'h42 == io_data_in[63:56] ? 8'h2c : _GEN_1601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1603 = 8'h43 == io_data_in[63:56] ? 8'h1a : _GEN_1602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1604 = 8'h44 == io_data_in[63:56] ? 8'h1b : _GEN_1603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1605 = 8'h45 == io_data_in[63:56] ? 8'h6e : _GEN_1604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1606 = 8'h46 == io_data_in[63:56] ? 8'h5a : _GEN_1605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1607 = 8'h47 == io_data_in[63:56] ? 8'ha0 : _GEN_1606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1608 = 8'h48 == io_data_in[63:56] ? 8'h52 : _GEN_1607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1609 = 8'h49 == io_data_in[63:56] ? 8'h3b : _GEN_1608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1610 = 8'h4a == io_data_in[63:56] ? 8'hd6 : _GEN_1609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1611 = 8'h4b == io_data_in[63:56] ? 8'hb3 : _GEN_1610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1612 = 8'h4c == io_data_in[63:56] ? 8'h29 : _GEN_1611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1613 = 8'h4d == io_data_in[63:56] ? 8'he3 : _GEN_1612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1614 = 8'h4e == io_data_in[63:56] ? 8'h2f : _GEN_1613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1615 = 8'h4f == io_data_in[63:56] ? 8'h84 : _GEN_1614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1616 = 8'h50 == io_data_in[63:56] ? 8'h53 : _GEN_1615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1617 = 8'h51 == io_data_in[63:56] ? 8'hd1 : _GEN_1616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1618 = 8'h52 == io_data_in[63:56] ? 8'h0 : _GEN_1617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1619 = 8'h53 == io_data_in[63:56] ? 8'hed : _GEN_1618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1620 = 8'h54 == io_data_in[63:56] ? 8'h20 : _GEN_1619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1621 = 8'h55 == io_data_in[63:56] ? 8'hfc : _GEN_1620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1622 = 8'h56 == io_data_in[63:56] ? 8'hb1 : _GEN_1621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1623 = 8'h57 == io_data_in[63:56] ? 8'h5b : _GEN_1622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1624 = 8'h58 == io_data_in[63:56] ? 8'h6a : _GEN_1623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1625 = 8'h59 == io_data_in[63:56] ? 8'hcb : _GEN_1624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1626 = 8'h5a == io_data_in[63:56] ? 8'hbe : _GEN_1625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1627 = 8'h5b == io_data_in[63:56] ? 8'h39 : _GEN_1626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1628 = 8'h5c == io_data_in[63:56] ? 8'h4a : _GEN_1627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1629 = 8'h5d == io_data_in[63:56] ? 8'h4c : _GEN_1628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1630 = 8'h5e == io_data_in[63:56] ? 8'h58 : _GEN_1629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1631 = 8'h5f == io_data_in[63:56] ? 8'hcf : _GEN_1630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1632 = 8'h60 == io_data_in[63:56] ? 8'hd0 : _GEN_1631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1633 = 8'h61 == io_data_in[63:56] ? 8'hef : _GEN_1632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1634 = 8'h62 == io_data_in[63:56] ? 8'haa : _GEN_1633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1635 = 8'h63 == io_data_in[63:56] ? 8'hfb : _GEN_1634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1636 = 8'h64 == io_data_in[63:56] ? 8'h43 : _GEN_1635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1637 = 8'h65 == io_data_in[63:56] ? 8'h4d : _GEN_1636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1638 = 8'h66 == io_data_in[63:56] ? 8'h33 : _GEN_1637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1639 = 8'h67 == io_data_in[63:56] ? 8'h85 : _GEN_1638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1640 = 8'h68 == io_data_in[63:56] ? 8'h45 : _GEN_1639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1641 = 8'h69 == io_data_in[63:56] ? 8'hf9 : _GEN_1640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1642 = 8'h6a == io_data_in[63:56] ? 8'h2 : _GEN_1641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1643 = 8'h6b == io_data_in[63:56] ? 8'h7f : _GEN_1642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1644 = 8'h6c == io_data_in[63:56] ? 8'h50 : _GEN_1643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1645 = 8'h6d == io_data_in[63:56] ? 8'h3c : _GEN_1644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1646 = 8'h6e == io_data_in[63:56] ? 8'h9f : _GEN_1645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1647 = 8'h6f == io_data_in[63:56] ? 8'ha8 : _GEN_1646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1648 = 8'h70 == io_data_in[63:56] ? 8'h51 : _GEN_1647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1649 = 8'h71 == io_data_in[63:56] ? 8'ha3 : _GEN_1648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1650 = 8'h72 == io_data_in[63:56] ? 8'h40 : _GEN_1649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1651 = 8'h73 == io_data_in[63:56] ? 8'h8f : _GEN_1650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1652 = 8'h74 == io_data_in[63:56] ? 8'h92 : _GEN_1651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1653 = 8'h75 == io_data_in[63:56] ? 8'h9d : _GEN_1652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1654 = 8'h76 == io_data_in[63:56] ? 8'h38 : _GEN_1653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1655 = 8'h77 == io_data_in[63:56] ? 8'hf5 : _GEN_1654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1656 = 8'h78 == io_data_in[63:56] ? 8'hbc : _GEN_1655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1657 = 8'h79 == io_data_in[63:56] ? 8'hb6 : _GEN_1656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1658 = 8'h7a == io_data_in[63:56] ? 8'hda : _GEN_1657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1659 = 8'h7b == io_data_in[63:56] ? 8'h21 : _GEN_1658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1660 = 8'h7c == io_data_in[63:56] ? 8'h10 : _GEN_1659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1661 = 8'h7d == io_data_in[63:56] ? 8'hff : _GEN_1660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1662 = 8'h7e == io_data_in[63:56] ? 8'hf3 : _GEN_1661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1663 = 8'h7f == io_data_in[63:56] ? 8'hd2 : _GEN_1662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1664 = 8'h80 == io_data_in[63:56] ? 8'hcd : _GEN_1663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1665 = 8'h81 == io_data_in[63:56] ? 8'hc : _GEN_1664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1666 = 8'h82 == io_data_in[63:56] ? 8'h13 : _GEN_1665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1667 = 8'h83 == io_data_in[63:56] ? 8'hec : _GEN_1666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1668 = 8'h84 == io_data_in[63:56] ? 8'h5f : _GEN_1667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1669 = 8'h85 == io_data_in[63:56] ? 8'h97 : _GEN_1668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1670 = 8'h86 == io_data_in[63:56] ? 8'h44 : _GEN_1669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1671 = 8'h87 == io_data_in[63:56] ? 8'h17 : _GEN_1670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1672 = 8'h88 == io_data_in[63:56] ? 8'hc4 : _GEN_1671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1673 = 8'h89 == io_data_in[63:56] ? 8'ha7 : _GEN_1672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1674 = 8'h8a == io_data_in[63:56] ? 8'h7e : _GEN_1673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1675 = 8'h8b == io_data_in[63:56] ? 8'h3d : _GEN_1674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1676 = 8'h8c == io_data_in[63:56] ? 8'h64 : _GEN_1675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1677 = 8'h8d == io_data_in[63:56] ? 8'h5d : _GEN_1676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1678 = 8'h8e == io_data_in[63:56] ? 8'h19 : _GEN_1677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1679 = 8'h8f == io_data_in[63:56] ? 8'h73 : _GEN_1678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1680 = 8'h90 == io_data_in[63:56] ? 8'h60 : _GEN_1679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1681 = 8'h91 == io_data_in[63:56] ? 8'h81 : _GEN_1680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1682 = 8'h92 == io_data_in[63:56] ? 8'h4f : _GEN_1681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1683 = 8'h93 == io_data_in[63:56] ? 8'hdc : _GEN_1682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1684 = 8'h94 == io_data_in[63:56] ? 8'h22 : _GEN_1683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1685 = 8'h95 == io_data_in[63:56] ? 8'h2a : _GEN_1684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1686 = 8'h96 == io_data_in[63:56] ? 8'h90 : _GEN_1685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1687 = 8'h97 == io_data_in[63:56] ? 8'h88 : _GEN_1686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1688 = 8'h98 == io_data_in[63:56] ? 8'h46 : _GEN_1687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1689 = 8'h99 == io_data_in[63:56] ? 8'hee : _GEN_1688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1690 = 8'h9a == io_data_in[63:56] ? 8'hb8 : _GEN_1689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1691 = 8'h9b == io_data_in[63:56] ? 8'h14 : _GEN_1690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1692 = 8'h9c == io_data_in[63:56] ? 8'hde : _GEN_1691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1693 = 8'h9d == io_data_in[63:56] ? 8'h5e : _GEN_1692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1694 = 8'h9e == io_data_in[63:56] ? 8'hb : _GEN_1693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1695 = 8'h9f == io_data_in[63:56] ? 8'hdb : _GEN_1694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1696 = 8'ha0 == io_data_in[63:56] ? 8'he0 : _GEN_1695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1697 = 8'ha1 == io_data_in[63:56] ? 8'h32 : _GEN_1696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1698 = 8'ha2 == io_data_in[63:56] ? 8'h3a : _GEN_1697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1699 = 8'ha3 == io_data_in[63:56] ? 8'ha : _GEN_1698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1700 = 8'ha4 == io_data_in[63:56] ? 8'h49 : _GEN_1699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1701 = 8'ha5 == io_data_in[63:56] ? 8'h6 : _GEN_1700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1702 = 8'ha6 == io_data_in[63:56] ? 8'h24 : _GEN_1701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1703 = 8'ha7 == io_data_in[63:56] ? 8'h5c : _GEN_1702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1704 = 8'ha8 == io_data_in[63:56] ? 8'hc2 : _GEN_1703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1705 = 8'ha9 == io_data_in[63:56] ? 8'hd3 : _GEN_1704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1706 = 8'haa == io_data_in[63:56] ? 8'hac : _GEN_1705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1707 = 8'hab == io_data_in[63:56] ? 8'h62 : _GEN_1706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1708 = 8'hac == io_data_in[63:56] ? 8'h91 : _GEN_1707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1709 = 8'had == io_data_in[63:56] ? 8'h95 : _GEN_1708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1710 = 8'hae == io_data_in[63:56] ? 8'he4 : _GEN_1709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1711 = 8'haf == io_data_in[63:56] ? 8'h79 : _GEN_1710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1712 = 8'hb0 == io_data_in[63:56] ? 8'he7 : _GEN_1711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1713 = 8'hb1 == io_data_in[63:56] ? 8'hc8 : _GEN_1712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1714 = 8'hb2 == io_data_in[63:56] ? 8'h37 : _GEN_1713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1715 = 8'hb3 == io_data_in[63:56] ? 8'h6d : _GEN_1714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1716 = 8'hb4 == io_data_in[63:56] ? 8'h8d : _GEN_1715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1717 = 8'hb5 == io_data_in[63:56] ? 8'hd5 : _GEN_1716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1718 = 8'hb6 == io_data_in[63:56] ? 8'h4e : _GEN_1717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1719 = 8'hb7 == io_data_in[63:56] ? 8'ha9 : _GEN_1718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1720 = 8'hb8 == io_data_in[63:56] ? 8'h6c : _GEN_1719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1721 = 8'hb9 == io_data_in[63:56] ? 8'h56 : _GEN_1720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1722 = 8'hba == io_data_in[63:56] ? 8'hf4 : _GEN_1721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1723 = 8'hbb == io_data_in[63:56] ? 8'hea : _GEN_1722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1724 = 8'hbc == io_data_in[63:56] ? 8'h65 : _GEN_1723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1725 = 8'hbd == io_data_in[63:56] ? 8'h7a : _GEN_1724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1726 = 8'hbe == io_data_in[63:56] ? 8'hae : _GEN_1725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1727 = 8'hbf == io_data_in[63:56] ? 8'h8 : _GEN_1726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1728 = 8'hc0 == io_data_in[63:56] ? 8'hba : _GEN_1727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1729 = 8'hc1 == io_data_in[63:56] ? 8'h78 : _GEN_1728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1730 = 8'hc2 == io_data_in[63:56] ? 8'h25 : _GEN_1729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1731 = 8'hc3 == io_data_in[63:56] ? 8'h2e : _GEN_1730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1732 = 8'hc4 == io_data_in[63:56] ? 8'h1c : _GEN_1731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1733 = 8'hc5 == io_data_in[63:56] ? 8'ha6 : _GEN_1732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1734 = 8'hc6 == io_data_in[63:56] ? 8'hb4 : _GEN_1733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1735 = 8'hc7 == io_data_in[63:56] ? 8'hc6 : _GEN_1734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1736 = 8'hc8 == io_data_in[63:56] ? 8'he8 : _GEN_1735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1737 = 8'hc9 == io_data_in[63:56] ? 8'hdd : _GEN_1736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1738 = 8'hca == io_data_in[63:56] ? 8'h74 : _GEN_1737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1739 = 8'hcb == io_data_in[63:56] ? 8'h1f : _GEN_1738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1740 = 8'hcc == io_data_in[63:56] ? 8'h4b : _GEN_1739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1741 = 8'hcd == io_data_in[63:56] ? 8'hbd : _GEN_1740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1742 = 8'hce == io_data_in[63:56] ? 8'h8b : _GEN_1741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1743 = 8'hcf == io_data_in[63:56] ? 8'h8a : _GEN_1742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1744 = 8'hd0 == io_data_in[63:56] ? 8'h70 : _GEN_1743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1745 = 8'hd1 == io_data_in[63:56] ? 8'h3e : _GEN_1744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1746 = 8'hd2 == io_data_in[63:56] ? 8'hb5 : _GEN_1745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1747 = 8'hd3 == io_data_in[63:56] ? 8'h66 : _GEN_1746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1748 = 8'hd4 == io_data_in[63:56] ? 8'h48 : _GEN_1747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1749 = 8'hd5 == io_data_in[63:56] ? 8'h3 : _GEN_1748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1750 = 8'hd6 == io_data_in[63:56] ? 8'hf6 : _GEN_1749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1751 = 8'hd7 == io_data_in[63:56] ? 8'he : _GEN_1750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1752 = 8'hd8 == io_data_in[63:56] ? 8'h61 : _GEN_1751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1753 = 8'hd9 == io_data_in[63:56] ? 8'h35 : _GEN_1752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1754 = 8'hda == io_data_in[63:56] ? 8'h57 : _GEN_1753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1755 = 8'hdb == io_data_in[63:56] ? 8'hb9 : _GEN_1754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1756 = 8'hdc == io_data_in[63:56] ? 8'h86 : _GEN_1755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1757 = 8'hdd == io_data_in[63:56] ? 8'hc1 : _GEN_1756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1758 = 8'hde == io_data_in[63:56] ? 8'h1d : _GEN_1757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1759 = 8'hdf == io_data_in[63:56] ? 8'h9e : _GEN_1758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1760 = 8'he0 == io_data_in[63:56] ? 8'he1 : _GEN_1759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1761 = 8'he1 == io_data_in[63:56] ? 8'hf8 : _GEN_1760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1762 = 8'he2 == io_data_in[63:56] ? 8'h98 : _GEN_1761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1763 = 8'he3 == io_data_in[63:56] ? 8'h11 : _GEN_1762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1764 = 8'he4 == io_data_in[63:56] ? 8'h69 : _GEN_1763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1765 = 8'he5 == io_data_in[63:56] ? 8'hd9 : _GEN_1764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1766 = 8'he6 == io_data_in[63:56] ? 8'h8e : _GEN_1765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1767 = 8'he7 == io_data_in[63:56] ? 8'h94 : _GEN_1766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1768 = 8'he8 == io_data_in[63:56] ? 8'h9b : _GEN_1767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1769 = 8'he9 == io_data_in[63:56] ? 8'h1e : _GEN_1768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1770 = 8'hea == io_data_in[63:56] ? 8'h87 : _GEN_1769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1771 = 8'heb == io_data_in[63:56] ? 8'he9 : _GEN_1770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1772 = 8'hec == io_data_in[63:56] ? 8'hce : _GEN_1771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1773 = 8'hed == io_data_in[63:56] ? 8'h55 : _GEN_1772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1774 = 8'hee == io_data_in[63:56] ? 8'h28 : _GEN_1773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1775 = 8'hef == io_data_in[63:56] ? 8'hdf : _GEN_1774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1776 = 8'hf0 == io_data_in[63:56] ? 8'h8c : _GEN_1775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1777 = 8'hf1 == io_data_in[63:56] ? 8'ha1 : _GEN_1776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1778 = 8'hf2 == io_data_in[63:56] ? 8'h89 : _GEN_1777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1779 = 8'hf3 == io_data_in[63:56] ? 8'hd : _GEN_1778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1780 = 8'hf4 == io_data_in[63:56] ? 8'hbf : _GEN_1779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1781 = 8'hf5 == io_data_in[63:56] ? 8'he6 : _GEN_1780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1782 = 8'hf6 == io_data_in[63:56] ? 8'h42 : _GEN_1781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1783 = 8'hf7 == io_data_in[63:56] ? 8'h68 : _GEN_1782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1784 = 8'hf8 == io_data_in[63:56] ? 8'h41 : _GEN_1783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1785 = 8'hf9 == io_data_in[63:56] ? 8'h99 : _GEN_1784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1786 = 8'hfa == io_data_in[63:56] ? 8'h2d : _GEN_1785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1787 = 8'hfb == io_data_in[63:56] ? 8'hf : _GEN_1786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1788 = 8'hfc == io_data_in[63:56] ? 8'hb0 : _GEN_1787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1789 = 8'hfd == io_data_in[63:56] ? 8'h54 : _GEN_1788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1790 = 8'hfe == io_data_in[63:56] ? 8'hbb : _GEN_1789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1791 = 8'hff == io_data_in[63:56] ? 8'h16 : _GEN_1790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1793 = 8'h1 == io_data_in[55:48] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1794 = 8'h2 == io_data_in[55:48] ? 8'h77 : _GEN_1793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1795 = 8'h3 == io_data_in[55:48] ? 8'h7b : _GEN_1794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1796 = 8'h4 == io_data_in[55:48] ? 8'hf2 : _GEN_1795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1797 = 8'h5 == io_data_in[55:48] ? 8'h6b : _GEN_1796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1798 = 8'h6 == io_data_in[55:48] ? 8'h6f : _GEN_1797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1799 = 8'h7 == io_data_in[55:48] ? 8'hc5 : _GEN_1798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1800 = 8'h8 == io_data_in[55:48] ? 8'h30 : _GEN_1799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1801 = 8'h9 == io_data_in[55:48] ? 8'h1 : _GEN_1800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1802 = 8'ha == io_data_in[55:48] ? 8'h67 : _GEN_1801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1803 = 8'hb == io_data_in[55:48] ? 8'h2b : _GEN_1802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1804 = 8'hc == io_data_in[55:48] ? 8'hfe : _GEN_1803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1805 = 8'hd == io_data_in[55:48] ? 8'hd7 : _GEN_1804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1806 = 8'he == io_data_in[55:48] ? 8'hab : _GEN_1805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1807 = 8'hf == io_data_in[55:48] ? 8'h76 : _GEN_1806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1808 = 8'h10 == io_data_in[55:48] ? 8'hca : _GEN_1807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1809 = 8'h11 == io_data_in[55:48] ? 8'h82 : _GEN_1808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1810 = 8'h12 == io_data_in[55:48] ? 8'hc9 : _GEN_1809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1811 = 8'h13 == io_data_in[55:48] ? 8'h7d : _GEN_1810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1812 = 8'h14 == io_data_in[55:48] ? 8'hfa : _GEN_1811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1813 = 8'h15 == io_data_in[55:48] ? 8'h59 : _GEN_1812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1814 = 8'h16 == io_data_in[55:48] ? 8'h47 : _GEN_1813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1815 = 8'h17 == io_data_in[55:48] ? 8'hf0 : _GEN_1814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1816 = 8'h18 == io_data_in[55:48] ? 8'had : _GEN_1815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1817 = 8'h19 == io_data_in[55:48] ? 8'hd4 : _GEN_1816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1818 = 8'h1a == io_data_in[55:48] ? 8'ha2 : _GEN_1817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1819 = 8'h1b == io_data_in[55:48] ? 8'haf : _GEN_1818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1820 = 8'h1c == io_data_in[55:48] ? 8'h9c : _GEN_1819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1821 = 8'h1d == io_data_in[55:48] ? 8'ha4 : _GEN_1820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1822 = 8'h1e == io_data_in[55:48] ? 8'h72 : _GEN_1821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1823 = 8'h1f == io_data_in[55:48] ? 8'hc0 : _GEN_1822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1824 = 8'h20 == io_data_in[55:48] ? 8'hb7 : _GEN_1823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1825 = 8'h21 == io_data_in[55:48] ? 8'hfd : _GEN_1824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1826 = 8'h22 == io_data_in[55:48] ? 8'h93 : _GEN_1825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1827 = 8'h23 == io_data_in[55:48] ? 8'h26 : _GEN_1826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1828 = 8'h24 == io_data_in[55:48] ? 8'h36 : _GEN_1827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1829 = 8'h25 == io_data_in[55:48] ? 8'h3f : _GEN_1828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1830 = 8'h26 == io_data_in[55:48] ? 8'hf7 : _GEN_1829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1831 = 8'h27 == io_data_in[55:48] ? 8'hcc : _GEN_1830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1832 = 8'h28 == io_data_in[55:48] ? 8'h34 : _GEN_1831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1833 = 8'h29 == io_data_in[55:48] ? 8'ha5 : _GEN_1832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1834 = 8'h2a == io_data_in[55:48] ? 8'he5 : _GEN_1833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1835 = 8'h2b == io_data_in[55:48] ? 8'hf1 : _GEN_1834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1836 = 8'h2c == io_data_in[55:48] ? 8'h71 : _GEN_1835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1837 = 8'h2d == io_data_in[55:48] ? 8'hd8 : _GEN_1836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1838 = 8'h2e == io_data_in[55:48] ? 8'h31 : _GEN_1837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1839 = 8'h2f == io_data_in[55:48] ? 8'h15 : _GEN_1838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1840 = 8'h30 == io_data_in[55:48] ? 8'h4 : _GEN_1839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1841 = 8'h31 == io_data_in[55:48] ? 8'hc7 : _GEN_1840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1842 = 8'h32 == io_data_in[55:48] ? 8'h23 : _GEN_1841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1843 = 8'h33 == io_data_in[55:48] ? 8'hc3 : _GEN_1842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1844 = 8'h34 == io_data_in[55:48] ? 8'h18 : _GEN_1843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1845 = 8'h35 == io_data_in[55:48] ? 8'h96 : _GEN_1844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1846 = 8'h36 == io_data_in[55:48] ? 8'h5 : _GEN_1845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1847 = 8'h37 == io_data_in[55:48] ? 8'h9a : _GEN_1846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1848 = 8'h38 == io_data_in[55:48] ? 8'h7 : _GEN_1847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1849 = 8'h39 == io_data_in[55:48] ? 8'h12 : _GEN_1848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1850 = 8'h3a == io_data_in[55:48] ? 8'h80 : _GEN_1849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1851 = 8'h3b == io_data_in[55:48] ? 8'he2 : _GEN_1850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1852 = 8'h3c == io_data_in[55:48] ? 8'heb : _GEN_1851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1853 = 8'h3d == io_data_in[55:48] ? 8'h27 : _GEN_1852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1854 = 8'h3e == io_data_in[55:48] ? 8'hb2 : _GEN_1853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1855 = 8'h3f == io_data_in[55:48] ? 8'h75 : _GEN_1854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1856 = 8'h40 == io_data_in[55:48] ? 8'h9 : _GEN_1855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1857 = 8'h41 == io_data_in[55:48] ? 8'h83 : _GEN_1856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1858 = 8'h42 == io_data_in[55:48] ? 8'h2c : _GEN_1857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1859 = 8'h43 == io_data_in[55:48] ? 8'h1a : _GEN_1858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1860 = 8'h44 == io_data_in[55:48] ? 8'h1b : _GEN_1859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1861 = 8'h45 == io_data_in[55:48] ? 8'h6e : _GEN_1860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1862 = 8'h46 == io_data_in[55:48] ? 8'h5a : _GEN_1861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1863 = 8'h47 == io_data_in[55:48] ? 8'ha0 : _GEN_1862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1864 = 8'h48 == io_data_in[55:48] ? 8'h52 : _GEN_1863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1865 = 8'h49 == io_data_in[55:48] ? 8'h3b : _GEN_1864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1866 = 8'h4a == io_data_in[55:48] ? 8'hd6 : _GEN_1865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1867 = 8'h4b == io_data_in[55:48] ? 8'hb3 : _GEN_1866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1868 = 8'h4c == io_data_in[55:48] ? 8'h29 : _GEN_1867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1869 = 8'h4d == io_data_in[55:48] ? 8'he3 : _GEN_1868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1870 = 8'h4e == io_data_in[55:48] ? 8'h2f : _GEN_1869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1871 = 8'h4f == io_data_in[55:48] ? 8'h84 : _GEN_1870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1872 = 8'h50 == io_data_in[55:48] ? 8'h53 : _GEN_1871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1873 = 8'h51 == io_data_in[55:48] ? 8'hd1 : _GEN_1872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1874 = 8'h52 == io_data_in[55:48] ? 8'h0 : _GEN_1873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1875 = 8'h53 == io_data_in[55:48] ? 8'hed : _GEN_1874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1876 = 8'h54 == io_data_in[55:48] ? 8'h20 : _GEN_1875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1877 = 8'h55 == io_data_in[55:48] ? 8'hfc : _GEN_1876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1878 = 8'h56 == io_data_in[55:48] ? 8'hb1 : _GEN_1877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1879 = 8'h57 == io_data_in[55:48] ? 8'h5b : _GEN_1878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1880 = 8'h58 == io_data_in[55:48] ? 8'h6a : _GEN_1879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1881 = 8'h59 == io_data_in[55:48] ? 8'hcb : _GEN_1880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1882 = 8'h5a == io_data_in[55:48] ? 8'hbe : _GEN_1881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1883 = 8'h5b == io_data_in[55:48] ? 8'h39 : _GEN_1882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1884 = 8'h5c == io_data_in[55:48] ? 8'h4a : _GEN_1883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1885 = 8'h5d == io_data_in[55:48] ? 8'h4c : _GEN_1884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1886 = 8'h5e == io_data_in[55:48] ? 8'h58 : _GEN_1885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1887 = 8'h5f == io_data_in[55:48] ? 8'hcf : _GEN_1886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1888 = 8'h60 == io_data_in[55:48] ? 8'hd0 : _GEN_1887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1889 = 8'h61 == io_data_in[55:48] ? 8'hef : _GEN_1888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1890 = 8'h62 == io_data_in[55:48] ? 8'haa : _GEN_1889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1891 = 8'h63 == io_data_in[55:48] ? 8'hfb : _GEN_1890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1892 = 8'h64 == io_data_in[55:48] ? 8'h43 : _GEN_1891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1893 = 8'h65 == io_data_in[55:48] ? 8'h4d : _GEN_1892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1894 = 8'h66 == io_data_in[55:48] ? 8'h33 : _GEN_1893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1895 = 8'h67 == io_data_in[55:48] ? 8'h85 : _GEN_1894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1896 = 8'h68 == io_data_in[55:48] ? 8'h45 : _GEN_1895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1897 = 8'h69 == io_data_in[55:48] ? 8'hf9 : _GEN_1896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1898 = 8'h6a == io_data_in[55:48] ? 8'h2 : _GEN_1897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1899 = 8'h6b == io_data_in[55:48] ? 8'h7f : _GEN_1898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1900 = 8'h6c == io_data_in[55:48] ? 8'h50 : _GEN_1899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1901 = 8'h6d == io_data_in[55:48] ? 8'h3c : _GEN_1900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1902 = 8'h6e == io_data_in[55:48] ? 8'h9f : _GEN_1901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1903 = 8'h6f == io_data_in[55:48] ? 8'ha8 : _GEN_1902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1904 = 8'h70 == io_data_in[55:48] ? 8'h51 : _GEN_1903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1905 = 8'h71 == io_data_in[55:48] ? 8'ha3 : _GEN_1904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1906 = 8'h72 == io_data_in[55:48] ? 8'h40 : _GEN_1905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1907 = 8'h73 == io_data_in[55:48] ? 8'h8f : _GEN_1906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1908 = 8'h74 == io_data_in[55:48] ? 8'h92 : _GEN_1907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1909 = 8'h75 == io_data_in[55:48] ? 8'h9d : _GEN_1908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1910 = 8'h76 == io_data_in[55:48] ? 8'h38 : _GEN_1909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1911 = 8'h77 == io_data_in[55:48] ? 8'hf5 : _GEN_1910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1912 = 8'h78 == io_data_in[55:48] ? 8'hbc : _GEN_1911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1913 = 8'h79 == io_data_in[55:48] ? 8'hb6 : _GEN_1912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1914 = 8'h7a == io_data_in[55:48] ? 8'hda : _GEN_1913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1915 = 8'h7b == io_data_in[55:48] ? 8'h21 : _GEN_1914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1916 = 8'h7c == io_data_in[55:48] ? 8'h10 : _GEN_1915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1917 = 8'h7d == io_data_in[55:48] ? 8'hff : _GEN_1916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1918 = 8'h7e == io_data_in[55:48] ? 8'hf3 : _GEN_1917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1919 = 8'h7f == io_data_in[55:48] ? 8'hd2 : _GEN_1918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1920 = 8'h80 == io_data_in[55:48] ? 8'hcd : _GEN_1919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1921 = 8'h81 == io_data_in[55:48] ? 8'hc : _GEN_1920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1922 = 8'h82 == io_data_in[55:48] ? 8'h13 : _GEN_1921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1923 = 8'h83 == io_data_in[55:48] ? 8'hec : _GEN_1922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1924 = 8'h84 == io_data_in[55:48] ? 8'h5f : _GEN_1923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1925 = 8'h85 == io_data_in[55:48] ? 8'h97 : _GEN_1924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1926 = 8'h86 == io_data_in[55:48] ? 8'h44 : _GEN_1925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1927 = 8'h87 == io_data_in[55:48] ? 8'h17 : _GEN_1926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1928 = 8'h88 == io_data_in[55:48] ? 8'hc4 : _GEN_1927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1929 = 8'h89 == io_data_in[55:48] ? 8'ha7 : _GEN_1928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1930 = 8'h8a == io_data_in[55:48] ? 8'h7e : _GEN_1929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1931 = 8'h8b == io_data_in[55:48] ? 8'h3d : _GEN_1930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1932 = 8'h8c == io_data_in[55:48] ? 8'h64 : _GEN_1931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1933 = 8'h8d == io_data_in[55:48] ? 8'h5d : _GEN_1932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1934 = 8'h8e == io_data_in[55:48] ? 8'h19 : _GEN_1933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1935 = 8'h8f == io_data_in[55:48] ? 8'h73 : _GEN_1934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1936 = 8'h90 == io_data_in[55:48] ? 8'h60 : _GEN_1935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1937 = 8'h91 == io_data_in[55:48] ? 8'h81 : _GEN_1936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1938 = 8'h92 == io_data_in[55:48] ? 8'h4f : _GEN_1937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1939 = 8'h93 == io_data_in[55:48] ? 8'hdc : _GEN_1938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1940 = 8'h94 == io_data_in[55:48] ? 8'h22 : _GEN_1939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1941 = 8'h95 == io_data_in[55:48] ? 8'h2a : _GEN_1940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1942 = 8'h96 == io_data_in[55:48] ? 8'h90 : _GEN_1941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1943 = 8'h97 == io_data_in[55:48] ? 8'h88 : _GEN_1942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1944 = 8'h98 == io_data_in[55:48] ? 8'h46 : _GEN_1943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1945 = 8'h99 == io_data_in[55:48] ? 8'hee : _GEN_1944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1946 = 8'h9a == io_data_in[55:48] ? 8'hb8 : _GEN_1945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1947 = 8'h9b == io_data_in[55:48] ? 8'h14 : _GEN_1946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1948 = 8'h9c == io_data_in[55:48] ? 8'hde : _GEN_1947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1949 = 8'h9d == io_data_in[55:48] ? 8'h5e : _GEN_1948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1950 = 8'h9e == io_data_in[55:48] ? 8'hb : _GEN_1949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1951 = 8'h9f == io_data_in[55:48] ? 8'hdb : _GEN_1950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1952 = 8'ha0 == io_data_in[55:48] ? 8'he0 : _GEN_1951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1953 = 8'ha1 == io_data_in[55:48] ? 8'h32 : _GEN_1952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1954 = 8'ha2 == io_data_in[55:48] ? 8'h3a : _GEN_1953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1955 = 8'ha3 == io_data_in[55:48] ? 8'ha : _GEN_1954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1956 = 8'ha4 == io_data_in[55:48] ? 8'h49 : _GEN_1955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1957 = 8'ha5 == io_data_in[55:48] ? 8'h6 : _GEN_1956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1958 = 8'ha6 == io_data_in[55:48] ? 8'h24 : _GEN_1957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1959 = 8'ha7 == io_data_in[55:48] ? 8'h5c : _GEN_1958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1960 = 8'ha8 == io_data_in[55:48] ? 8'hc2 : _GEN_1959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1961 = 8'ha9 == io_data_in[55:48] ? 8'hd3 : _GEN_1960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1962 = 8'haa == io_data_in[55:48] ? 8'hac : _GEN_1961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1963 = 8'hab == io_data_in[55:48] ? 8'h62 : _GEN_1962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1964 = 8'hac == io_data_in[55:48] ? 8'h91 : _GEN_1963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1965 = 8'had == io_data_in[55:48] ? 8'h95 : _GEN_1964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1966 = 8'hae == io_data_in[55:48] ? 8'he4 : _GEN_1965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1967 = 8'haf == io_data_in[55:48] ? 8'h79 : _GEN_1966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1968 = 8'hb0 == io_data_in[55:48] ? 8'he7 : _GEN_1967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1969 = 8'hb1 == io_data_in[55:48] ? 8'hc8 : _GEN_1968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1970 = 8'hb2 == io_data_in[55:48] ? 8'h37 : _GEN_1969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1971 = 8'hb3 == io_data_in[55:48] ? 8'h6d : _GEN_1970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1972 = 8'hb4 == io_data_in[55:48] ? 8'h8d : _GEN_1971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1973 = 8'hb5 == io_data_in[55:48] ? 8'hd5 : _GEN_1972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1974 = 8'hb6 == io_data_in[55:48] ? 8'h4e : _GEN_1973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1975 = 8'hb7 == io_data_in[55:48] ? 8'ha9 : _GEN_1974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1976 = 8'hb8 == io_data_in[55:48] ? 8'h6c : _GEN_1975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1977 = 8'hb9 == io_data_in[55:48] ? 8'h56 : _GEN_1976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1978 = 8'hba == io_data_in[55:48] ? 8'hf4 : _GEN_1977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1979 = 8'hbb == io_data_in[55:48] ? 8'hea : _GEN_1978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1980 = 8'hbc == io_data_in[55:48] ? 8'h65 : _GEN_1979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1981 = 8'hbd == io_data_in[55:48] ? 8'h7a : _GEN_1980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1982 = 8'hbe == io_data_in[55:48] ? 8'hae : _GEN_1981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1983 = 8'hbf == io_data_in[55:48] ? 8'h8 : _GEN_1982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1984 = 8'hc0 == io_data_in[55:48] ? 8'hba : _GEN_1983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1985 = 8'hc1 == io_data_in[55:48] ? 8'h78 : _GEN_1984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1986 = 8'hc2 == io_data_in[55:48] ? 8'h25 : _GEN_1985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1987 = 8'hc3 == io_data_in[55:48] ? 8'h2e : _GEN_1986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1988 = 8'hc4 == io_data_in[55:48] ? 8'h1c : _GEN_1987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1989 = 8'hc5 == io_data_in[55:48] ? 8'ha6 : _GEN_1988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1990 = 8'hc6 == io_data_in[55:48] ? 8'hb4 : _GEN_1989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1991 = 8'hc7 == io_data_in[55:48] ? 8'hc6 : _GEN_1990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1992 = 8'hc8 == io_data_in[55:48] ? 8'he8 : _GEN_1991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1993 = 8'hc9 == io_data_in[55:48] ? 8'hdd : _GEN_1992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1994 = 8'hca == io_data_in[55:48] ? 8'h74 : _GEN_1993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1995 = 8'hcb == io_data_in[55:48] ? 8'h1f : _GEN_1994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1996 = 8'hcc == io_data_in[55:48] ? 8'h4b : _GEN_1995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1997 = 8'hcd == io_data_in[55:48] ? 8'hbd : _GEN_1996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1998 = 8'hce == io_data_in[55:48] ? 8'h8b : _GEN_1997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1999 = 8'hcf == io_data_in[55:48] ? 8'h8a : _GEN_1998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2000 = 8'hd0 == io_data_in[55:48] ? 8'h70 : _GEN_1999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2001 = 8'hd1 == io_data_in[55:48] ? 8'h3e : _GEN_2000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2002 = 8'hd2 == io_data_in[55:48] ? 8'hb5 : _GEN_2001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2003 = 8'hd3 == io_data_in[55:48] ? 8'h66 : _GEN_2002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2004 = 8'hd4 == io_data_in[55:48] ? 8'h48 : _GEN_2003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2005 = 8'hd5 == io_data_in[55:48] ? 8'h3 : _GEN_2004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2006 = 8'hd6 == io_data_in[55:48] ? 8'hf6 : _GEN_2005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2007 = 8'hd7 == io_data_in[55:48] ? 8'he : _GEN_2006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2008 = 8'hd8 == io_data_in[55:48] ? 8'h61 : _GEN_2007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2009 = 8'hd9 == io_data_in[55:48] ? 8'h35 : _GEN_2008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2010 = 8'hda == io_data_in[55:48] ? 8'h57 : _GEN_2009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2011 = 8'hdb == io_data_in[55:48] ? 8'hb9 : _GEN_2010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2012 = 8'hdc == io_data_in[55:48] ? 8'h86 : _GEN_2011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2013 = 8'hdd == io_data_in[55:48] ? 8'hc1 : _GEN_2012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2014 = 8'hde == io_data_in[55:48] ? 8'h1d : _GEN_2013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2015 = 8'hdf == io_data_in[55:48] ? 8'h9e : _GEN_2014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2016 = 8'he0 == io_data_in[55:48] ? 8'he1 : _GEN_2015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2017 = 8'he1 == io_data_in[55:48] ? 8'hf8 : _GEN_2016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2018 = 8'he2 == io_data_in[55:48] ? 8'h98 : _GEN_2017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2019 = 8'he3 == io_data_in[55:48] ? 8'h11 : _GEN_2018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2020 = 8'he4 == io_data_in[55:48] ? 8'h69 : _GEN_2019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2021 = 8'he5 == io_data_in[55:48] ? 8'hd9 : _GEN_2020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2022 = 8'he6 == io_data_in[55:48] ? 8'h8e : _GEN_2021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2023 = 8'he7 == io_data_in[55:48] ? 8'h94 : _GEN_2022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2024 = 8'he8 == io_data_in[55:48] ? 8'h9b : _GEN_2023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2025 = 8'he9 == io_data_in[55:48] ? 8'h1e : _GEN_2024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2026 = 8'hea == io_data_in[55:48] ? 8'h87 : _GEN_2025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2027 = 8'heb == io_data_in[55:48] ? 8'he9 : _GEN_2026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2028 = 8'hec == io_data_in[55:48] ? 8'hce : _GEN_2027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2029 = 8'hed == io_data_in[55:48] ? 8'h55 : _GEN_2028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2030 = 8'hee == io_data_in[55:48] ? 8'h28 : _GEN_2029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2031 = 8'hef == io_data_in[55:48] ? 8'hdf : _GEN_2030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2032 = 8'hf0 == io_data_in[55:48] ? 8'h8c : _GEN_2031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2033 = 8'hf1 == io_data_in[55:48] ? 8'ha1 : _GEN_2032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2034 = 8'hf2 == io_data_in[55:48] ? 8'h89 : _GEN_2033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2035 = 8'hf3 == io_data_in[55:48] ? 8'hd : _GEN_2034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2036 = 8'hf4 == io_data_in[55:48] ? 8'hbf : _GEN_2035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2037 = 8'hf5 == io_data_in[55:48] ? 8'he6 : _GEN_2036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2038 = 8'hf6 == io_data_in[55:48] ? 8'h42 : _GEN_2037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2039 = 8'hf7 == io_data_in[55:48] ? 8'h68 : _GEN_2038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2040 = 8'hf8 == io_data_in[55:48] ? 8'h41 : _GEN_2039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2041 = 8'hf9 == io_data_in[55:48] ? 8'h99 : _GEN_2040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2042 = 8'hfa == io_data_in[55:48] ? 8'h2d : _GEN_2041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2043 = 8'hfb == io_data_in[55:48] ? 8'hf : _GEN_2042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2044 = 8'hfc == io_data_in[55:48] ? 8'hb0 : _GEN_2043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2045 = 8'hfd == io_data_in[55:48] ? 8'h54 : _GEN_2044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2046 = 8'hfe == io_data_in[55:48] ? 8'hbb : _GEN_2045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2047 = 8'hff == io_data_in[55:48] ? 8'h16 : _GEN_2046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [63:0] io_data_out_lo = {_GEN_1791,_GEN_2047,_GEN_1279,_GEN_1535,_GEN_767,_GEN_1023,_GEN_255,_GEN_511}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_2049 = 8'h1 == io_data_in[79:72] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2050 = 8'h2 == io_data_in[79:72] ? 8'h77 : _GEN_2049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2051 = 8'h3 == io_data_in[79:72] ? 8'h7b : _GEN_2050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2052 = 8'h4 == io_data_in[79:72] ? 8'hf2 : _GEN_2051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2053 = 8'h5 == io_data_in[79:72] ? 8'h6b : _GEN_2052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2054 = 8'h6 == io_data_in[79:72] ? 8'h6f : _GEN_2053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2055 = 8'h7 == io_data_in[79:72] ? 8'hc5 : _GEN_2054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2056 = 8'h8 == io_data_in[79:72] ? 8'h30 : _GEN_2055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2057 = 8'h9 == io_data_in[79:72] ? 8'h1 : _GEN_2056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2058 = 8'ha == io_data_in[79:72] ? 8'h67 : _GEN_2057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2059 = 8'hb == io_data_in[79:72] ? 8'h2b : _GEN_2058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2060 = 8'hc == io_data_in[79:72] ? 8'hfe : _GEN_2059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2061 = 8'hd == io_data_in[79:72] ? 8'hd7 : _GEN_2060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2062 = 8'he == io_data_in[79:72] ? 8'hab : _GEN_2061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2063 = 8'hf == io_data_in[79:72] ? 8'h76 : _GEN_2062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2064 = 8'h10 == io_data_in[79:72] ? 8'hca : _GEN_2063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2065 = 8'h11 == io_data_in[79:72] ? 8'h82 : _GEN_2064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2066 = 8'h12 == io_data_in[79:72] ? 8'hc9 : _GEN_2065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2067 = 8'h13 == io_data_in[79:72] ? 8'h7d : _GEN_2066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2068 = 8'h14 == io_data_in[79:72] ? 8'hfa : _GEN_2067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2069 = 8'h15 == io_data_in[79:72] ? 8'h59 : _GEN_2068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2070 = 8'h16 == io_data_in[79:72] ? 8'h47 : _GEN_2069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2071 = 8'h17 == io_data_in[79:72] ? 8'hf0 : _GEN_2070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2072 = 8'h18 == io_data_in[79:72] ? 8'had : _GEN_2071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2073 = 8'h19 == io_data_in[79:72] ? 8'hd4 : _GEN_2072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2074 = 8'h1a == io_data_in[79:72] ? 8'ha2 : _GEN_2073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2075 = 8'h1b == io_data_in[79:72] ? 8'haf : _GEN_2074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2076 = 8'h1c == io_data_in[79:72] ? 8'h9c : _GEN_2075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2077 = 8'h1d == io_data_in[79:72] ? 8'ha4 : _GEN_2076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2078 = 8'h1e == io_data_in[79:72] ? 8'h72 : _GEN_2077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2079 = 8'h1f == io_data_in[79:72] ? 8'hc0 : _GEN_2078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2080 = 8'h20 == io_data_in[79:72] ? 8'hb7 : _GEN_2079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2081 = 8'h21 == io_data_in[79:72] ? 8'hfd : _GEN_2080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2082 = 8'h22 == io_data_in[79:72] ? 8'h93 : _GEN_2081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2083 = 8'h23 == io_data_in[79:72] ? 8'h26 : _GEN_2082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2084 = 8'h24 == io_data_in[79:72] ? 8'h36 : _GEN_2083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2085 = 8'h25 == io_data_in[79:72] ? 8'h3f : _GEN_2084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2086 = 8'h26 == io_data_in[79:72] ? 8'hf7 : _GEN_2085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2087 = 8'h27 == io_data_in[79:72] ? 8'hcc : _GEN_2086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2088 = 8'h28 == io_data_in[79:72] ? 8'h34 : _GEN_2087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2089 = 8'h29 == io_data_in[79:72] ? 8'ha5 : _GEN_2088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2090 = 8'h2a == io_data_in[79:72] ? 8'he5 : _GEN_2089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2091 = 8'h2b == io_data_in[79:72] ? 8'hf1 : _GEN_2090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2092 = 8'h2c == io_data_in[79:72] ? 8'h71 : _GEN_2091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2093 = 8'h2d == io_data_in[79:72] ? 8'hd8 : _GEN_2092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2094 = 8'h2e == io_data_in[79:72] ? 8'h31 : _GEN_2093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2095 = 8'h2f == io_data_in[79:72] ? 8'h15 : _GEN_2094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2096 = 8'h30 == io_data_in[79:72] ? 8'h4 : _GEN_2095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2097 = 8'h31 == io_data_in[79:72] ? 8'hc7 : _GEN_2096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2098 = 8'h32 == io_data_in[79:72] ? 8'h23 : _GEN_2097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2099 = 8'h33 == io_data_in[79:72] ? 8'hc3 : _GEN_2098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2100 = 8'h34 == io_data_in[79:72] ? 8'h18 : _GEN_2099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2101 = 8'h35 == io_data_in[79:72] ? 8'h96 : _GEN_2100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2102 = 8'h36 == io_data_in[79:72] ? 8'h5 : _GEN_2101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2103 = 8'h37 == io_data_in[79:72] ? 8'h9a : _GEN_2102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2104 = 8'h38 == io_data_in[79:72] ? 8'h7 : _GEN_2103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2105 = 8'h39 == io_data_in[79:72] ? 8'h12 : _GEN_2104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2106 = 8'h3a == io_data_in[79:72] ? 8'h80 : _GEN_2105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2107 = 8'h3b == io_data_in[79:72] ? 8'he2 : _GEN_2106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2108 = 8'h3c == io_data_in[79:72] ? 8'heb : _GEN_2107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2109 = 8'h3d == io_data_in[79:72] ? 8'h27 : _GEN_2108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2110 = 8'h3e == io_data_in[79:72] ? 8'hb2 : _GEN_2109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2111 = 8'h3f == io_data_in[79:72] ? 8'h75 : _GEN_2110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2112 = 8'h40 == io_data_in[79:72] ? 8'h9 : _GEN_2111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2113 = 8'h41 == io_data_in[79:72] ? 8'h83 : _GEN_2112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2114 = 8'h42 == io_data_in[79:72] ? 8'h2c : _GEN_2113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2115 = 8'h43 == io_data_in[79:72] ? 8'h1a : _GEN_2114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2116 = 8'h44 == io_data_in[79:72] ? 8'h1b : _GEN_2115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2117 = 8'h45 == io_data_in[79:72] ? 8'h6e : _GEN_2116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2118 = 8'h46 == io_data_in[79:72] ? 8'h5a : _GEN_2117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2119 = 8'h47 == io_data_in[79:72] ? 8'ha0 : _GEN_2118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2120 = 8'h48 == io_data_in[79:72] ? 8'h52 : _GEN_2119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2121 = 8'h49 == io_data_in[79:72] ? 8'h3b : _GEN_2120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2122 = 8'h4a == io_data_in[79:72] ? 8'hd6 : _GEN_2121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2123 = 8'h4b == io_data_in[79:72] ? 8'hb3 : _GEN_2122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2124 = 8'h4c == io_data_in[79:72] ? 8'h29 : _GEN_2123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2125 = 8'h4d == io_data_in[79:72] ? 8'he3 : _GEN_2124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2126 = 8'h4e == io_data_in[79:72] ? 8'h2f : _GEN_2125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2127 = 8'h4f == io_data_in[79:72] ? 8'h84 : _GEN_2126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2128 = 8'h50 == io_data_in[79:72] ? 8'h53 : _GEN_2127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2129 = 8'h51 == io_data_in[79:72] ? 8'hd1 : _GEN_2128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2130 = 8'h52 == io_data_in[79:72] ? 8'h0 : _GEN_2129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2131 = 8'h53 == io_data_in[79:72] ? 8'hed : _GEN_2130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2132 = 8'h54 == io_data_in[79:72] ? 8'h20 : _GEN_2131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2133 = 8'h55 == io_data_in[79:72] ? 8'hfc : _GEN_2132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2134 = 8'h56 == io_data_in[79:72] ? 8'hb1 : _GEN_2133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2135 = 8'h57 == io_data_in[79:72] ? 8'h5b : _GEN_2134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2136 = 8'h58 == io_data_in[79:72] ? 8'h6a : _GEN_2135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2137 = 8'h59 == io_data_in[79:72] ? 8'hcb : _GEN_2136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2138 = 8'h5a == io_data_in[79:72] ? 8'hbe : _GEN_2137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2139 = 8'h5b == io_data_in[79:72] ? 8'h39 : _GEN_2138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2140 = 8'h5c == io_data_in[79:72] ? 8'h4a : _GEN_2139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2141 = 8'h5d == io_data_in[79:72] ? 8'h4c : _GEN_2140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2142 = 8'h5e == io_data_in[79:72] ? 8'h58 : _GEN_2141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2143 = 8'h5f == io_data_in[79:72] ? 8'hcf : _GEN_2142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2144 = 8'h60 == io_data_in[79:72] ? 8'hd0 : _GEN_2143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2145 = 8'h61 == io_data_in[79:72] ? 8'hef : _GEN_2144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2146 = 8'h62 == io_data_in[79:72] ? 8'haa : _GEN_2145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2147 = 8'h63 == io_data_in[79:72] ? 8'hfb : _GEN_2146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2148 = 8'h64 == io_data_in[79:72] ? 8'h43 : _GEN_2147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2149 = 8'h65 == io_data_in[79:72] ? 8'h4d : _GEN_2148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2150 = 8'h66 == io_data_in[79:72] ? 8'h33 : _GEN_2149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2151 = 8'h67 == io_data_in[79:72] ? 8'h85 : _GEN_2150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2152 = 8'h68 == io_data_in[79:72] ? 8'h45 : _GEN_2151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2153 = 8'h69 == io_data_in[79:72] ? 8'hf9 : _GEN_2152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2154 = 8'h6a == io_data_in[79:72] ? 8'h2 : _GEN_2153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2155 = 8'h6b == io_data_in[79:72] ? 8'h7f : _GEN_2154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2156 = 8'h6c == io_data_in[79:72] ? 8'h50 : _GEN_2155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2157 = 8'h6d == io_data_in[79:72] ? 8'h3c : _GEN_2156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2158 = 8'h6e == io_data_in[79:72] ? 8'h9f : _GEN_2157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2159 = 8'h6f == io_data_in[79:72] ? 8'ha8 : _GEN_2158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2160 = 8'h70 == io_data_in[79:72] ? 8'h51 : _GEN_2159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2161 = 8'h71 == io_data_in[79:72] ? 8'ha3 : _GEN_2160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2162 = 8'h72 == io_data_in[79:72] ? 8'h40 : _GEN_2161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2163 = 8'h73 == io_data_in[79:72] ? 8'h8f : _GEN_2162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2164 = 8'h74 == io_data_in[79:72] ? 8'h92 : _GEN_2163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2165 = 8'h75 == io_data_in[79:72] ? 8'h9d : _GEN_2164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2166 = 8'h76 == io_data_in[79:72] ? 8'h38 : _GEN_2165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2167 = 8'h77 == io_data_in[79:72] ? 8'hf5 : _GEN_2166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2168 = 8'h78 == io_data_in[79:72] ? 8'hbc : _GEN_2167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2169 = 8'h79 == io_data_in[79:72] ? 8'hb6 : _GEN_2168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2170 = 8'h7a == io_data_in[79:72] ? 8'hda : _GEN_2169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2171 = 8'h7b == io_data_in[79:72] ? 8'h21 : _GEN_2170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2172 = 8'h7c == io_data_in[79:72] ? 8'h10 : _GEN_2171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2173 = 8'h7d == io_data_in[79:72] ? 8'hff : _GEN_2172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2174 = 8'h7e == io_data_in[79:72] ? 8'hf3 : _GEN_2173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2175 = 8'h7f == io_data_in[79:72] ? 8'hd2 : _GEN_2174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2176 = 8'h80 == io_data_in[79:72] ? 8'hcd : _GEN_2175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2177 = 8'h81 == io_data_in[79:72] ? 8'hc : _GEN_2176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2178 = 8'h82 == io_data_in[79:72] ? 8'h13 : _GEN_2177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2179 = 8'h83 == io_data_in[79:72] ? 8'hec : _GEN_2178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2180 = 8'h84 == io_data_in[79:72] ? 8'h5f : _GEN_2179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2181 = 8'h85 == io_data_in[79:72] ? 8'h97 : _GEN_2180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2182 = 8'h86 == io_data_in[79:72] ? 8'h44 : _GEN_2181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2183 = 8'h87 == io_data_in[79:72] ? 8'h17 : _GEN_2182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2184 = 8'h88 == io_data_in[79:72] ? 8'hc4 : _GEN_2183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2185 = 8'h89 == io_data_in[79:72] ? 8'ha7 : _GEN_2184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2186 = 8'h8a == io_data_in[79:72] ? 8'h7e : _GEN_2185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2187 = 8'h8b == io_data_in[79:72] ? 8'h3d : _GEN_2186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2188 = 8'h8c == io_data_in[79:72] ? 8'h64 : _GEN_2187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2189 = 8'h8d == io_data_in[79:72] ? 8'h5d : _GEN_2188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2190 = 8'h8e == io_data_in[79:72] ? 8'h19 : _GEN_2189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2191 = 8'h8f == io_data_in[79:72] ? 8'h73 : _GEN_2190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2192 = 8'h90 == io_data_in[79:72] ? 8'h60 : _GEN_2191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2193 = 8'h91 == io_data_in[79:72] ? 8'h81 : _GEN_2192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2194 = 8'h92 == io_data_in[79:72] ? 8'h4f : _GEN_2193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2195 = 8'h93 == io_data_in[79:72] ? 8'hdc : _GEN_2194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2196 = 8'h94 == io_data_in[79:72] ? 8'h22 : _GEN_2195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2197 = 8'h95 == io_data_in[79:72] ? 8'h2a : _GEN_2196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2198 = 8'h96 == io_data_in[79:72] ? 8'h90 : _GEN_2197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2199 = 8'h97 == io_data_in[79:72] ? 8'h88 : _GEN_2198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2200 = 8'h98 == io_data_in[79:72] ? 8'h46 : _GEN_2199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2201 = 8'h99 == io_data_in[79:72] ? 8'hee : _GEN_2200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2202 = 8'h9a == io_data_in[79:72] ? 8'hb8 : _GEN_2201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2203 = 8'h9b == io_data_in[79:72] ? 8'h14 : _GEN_2202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2204 = 8'h9c == io_data_in[79:72] ? 8'hde : _GEN_2203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2205 = 8'h9d == io_data_in[79:72] ? 8'h5e : _GEN_2204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2206 = 8'h9e == io_data_in[79:72] ? 8'hb : _GEN_2205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2207 = 8'h9f == io_data_in[79:72] ? 8'hdb : _GEN_2206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2208 = 8'ha0 == io_data_in[79:72] ? 8'he0 : _GEN_2207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2209 = 8'ha1 == io_data_in[79:72] ? 8'h32 : _GEN_2208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2210 = 8'ha2 == io_data_in[79:72] ? 8'h3a : _GEN_2209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2211 = 8'ha3 == io_data_in[79:72] ? 8'ha : _GEN_2210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2212 = 8'ha4 == io_data_in[79:72] ? 8'h49 : _GEN_2211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2213 = 8'ha5 == io_data_in[79:72] ? 8'h6 : _GEN_2212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2214 = 8'ha6 == io_data_in[79:72] ? 8'h24 : _GEN_2213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2215 = 8'ha7 == io_data_in[79:72] ? 8'h5c : _GEN_2214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2216 = 8'ha8 == io_data_in[79:72] ? 8'hc2 : _GEN_2215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2217 = 8'ha9 == io_data_in[79:72] ? 8'hd3 : _GEN_2216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2218 = 8'haa == io_data_in[79:72] ? 8'hac : _GEN_2217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2219 = 8'hab == io_data_in[79:72] ? 8'h62 : _GEN_2218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2220 = 8'hac == io_data_in[79:72] ? 8'h91 : _GEN_2219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2221 = 8'had == io_data_in[79:72] ? 8'h95 : _GEN_2220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2222 = 8'hae == io_data_in[79:72] ? 8'he4 : _GEN_2221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2223 = 8'haf == io_data_in[79:72] ? 8'h79 : _GEN_2222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2224 = 8'hb0 == io_data_in[79:72] ? 8'he7 : _GEN_2223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2225 = 8'hb1 == io_data_in[79:72] ? 8'hc8 : _GEN_2224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2226 = 8'hb2 == io_data_in[79:72] ? 8'h37 : _GEN_2225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2227 = 8'hb3 == io_data_in[79:72] ? 8'h6d : _GEN_2226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2228 = 8'hb4 == io_data_in[79:72] ? 8'h8d : _GEN_2227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2229 = 8'hb5 == io_data_in[79:72] ? 8'hd5 : _GEN_2228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2230 = 8'hb6 == io_data_in[79:72] ? 8'h4e : _GEN_2229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2231 = 8'hb7 == io_data_in[79:72] ? 8'ha9 : _GEN_2230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2232 = 8'hb8 == io_data_in[79:72] ? 8'h6c : _GEN_2231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2233 = 8'hb9 == io_data_in[79:72] ? 8'h56 : _GEN_2232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2234 = 8'hba == io_data_in[79:72] ? 8'hf4 : _GEN_2233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2235 = 8'hbb == io_data_in[79:72] ? 8'hea : _GEN_2234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2236 = 8'hbc == io_data_in[79:72] ? 8'h65 : _GEN_2235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2237 = 8'hbd == io_data_in[79:72] ? 8'h7a : _GEN_2236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2238 = 8'hbe == io_data_in[79:72] ? 8'hae : _GEN_2237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2239 = 8'hbf == io_data_in[79:72] ? 8'h8 : _GEN_2238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2240 = 8'hc0 == io_data_in[79:72] ? 8'hba : _GEN_2239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2241 = 8'hc1 == io_data_in[79:72] ? 8'h78 : _GEN_2240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2242 = 8'hc2 == io_data_in[79:72] ? 8'h25 : _GEN_2241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2243 = 8'hc3 == io_data_in[79:72] ? 8'h2e : _GEN_2242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2244 = 8'hc4 == io_data_in[79:72] ? 8'h1c : _GEN_2243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2245 = 8'hc5 == io_data_in[79:72] ? 8'ha6 : _GEN_2244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2246 = 8'hc6 == io_data_in[79:72] ? 8'hb4 : _GEN_2245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2247 = 8'hc7 == io_data_in[79:72] ? 8'hc6 : _GEN_2246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2248 = 8'hc8 == io_data_in[79:72] ? 8'he8 : _GEN_2247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2249 = 8'hc9 == io_data_in[79:72] ? 8'hdd : _GEN_2248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2250 = 8'hca == io_data_in[79:72] ? 8'h74 : _GEN_2249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2251 = 8'hcb == io_data_in[79:72] ? 8'h1f : _GEN_2250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2252 = 8'hcc == io_data_in[79:72] ? 8'h4b : _GEN_2251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2253 = 8'hcd == io_data_in[79:72] ? 8'hbd : _GEN_2252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2254 = 8'hce == io_data_in[79:72] ? 8'h8b : _GEN_2253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2255 = 8'hcf == io_data_in[79:72] ? 8'h8a : _GEN_2254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2256 = 8'hd0 == io_data_in[79:72] ? 8'h70 : _GEN_2255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2257 = 8'hd1 == io_data_in[79:72] ? 8'h3e : _GEN_2256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2258 = 8'hd2 == io_data_in[79:72] ? 8'hb5 : _GEN_2257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2259 = 8'hd3 == io_data_in[79:72] ? 8'h66 : _GEN_2258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2260 = 8'hd4 == io_data_in[79:72] ? 8'h48 : _GEN_2259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2261 = 8'hd5 == io_data_in[79:72] ? 8'h3 : _GEN_2260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2262 = 8'hd6 == io_data_in[79:72] ? 8'hf6 : _GEN_2261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2263 = 8'hd7 == io_data_in[79:72] ? 8'he : _GEN_2262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2264 = 8'hd8 == io_data_in[79:72] ? 8'h61 : _GEN_2263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2265 = 8'hd9 == io_data_in[79:72] ? 8'h35 : _GEN_2264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2266 = 8'hda == io_data_in[79:72] ? 8'h57 : _GEN_2265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2267 = 8'hdb == io_data_in[79:72] ? 8'hb9 : _GEN_2266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2268 = 8'hdc == io_data_in[79:72] ? 8'h86 : _GEN_2267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2269 = 8'hdd == io_data_in[79:72] ? 8'hc1 : _GEN_2268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2270 = 8'hde == io_data_in[79:72] ? 8'h1d : _GEN_2269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2271 = 8'hdf == io_data_in[79:72] ? 8'h9e : _GEN_2270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2272 = 8'he0 == io_data_in[79:72] ? 8'he1 : _GEN_2271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2273 = 8'he1 == io_data_in[79:72] ? 8'hf8 : _GEN_2272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2274 = 8'he2 == io_data_in[79:72] ? 8'h98 : _GEN_2273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2275 = 8'he3 == io_data_in[79:72] ? 8'h11 : _GEN_2274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2276 = 8'he4 == io_data_in[79:72] ? 8'h69 : _GEN_2275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2277 = 8'he5 == io_data_in[79:72] ? 8'hd9 : _GEN_2276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2278 = 8'he6 == io_data_in[79:72] ? 8'h8e : _GEN_2277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2279 = 8'he7 == io_data_in[79:72] ? 8'h94 : _GEN_2278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2280 = 8'he8 == io_data_in[79:72] ? 8'h9b : _GEN_2279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2281 = 8'he9 == io_data_in[79:72] ? 8'h1e : _GEN_2280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2282 = 8'hea == io_data_in[79:72] ? 8'h87 : _GEN_2281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2283 = 8'heb == io_data_in[79:72] ? 8'he9 : _GEN_2282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2284 = 8'hec == io_data_in[79:72] ? 8'hce : _GEN_2283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2285 = 8'hed == io_data_in[79:72] ? 8'h55 : _GEN_2284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2286 = 8'hee == io_data_in[79:72] ? 8'h28 : _GEN_2285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2287 = 8'hef == io_data_in[79:72] ? 8'hdf : _GEN_2286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2288 = 8'hf0 == io_data_in[79:72] ? 8'h8c : _GEN_2287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2289 = 8'hf1 == io_data_in[79:72] ? 8'ha1 : _GEN_2288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2290 = 8'hf2 == io_data_in[79:72] ? 8'h89 : _GEN_2289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2291 = 8'hf3 == io_data_in[79:72] ? 8'hd : _GEN_2290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2292 = 8'hf4 == io_data_in[79:72] ? 8'hbf : _GEN_2291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2293 = 8'hf5 == io_data_in[79:72] ? 8'he6 : _GEN_2292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2294 = 8'hf6 == io_data_in[79:72] ? 8'h42 : _GEN_2293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2295 = 8'hf7 == io_data_in[79:72] ? 8'h68 : _GEN_2294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2296 = 8'hf8 == io_data_in[79:72] ? 8'h41 : _GEN_2295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2297 = 8'hf9 == io_data_in[79:72] ? 8'h99 : _GEN_2296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2298 = 8'hfa == io_data_in[79:72] ? 8'h2d : _GEN_2297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2299 = 8'hfb == io_data_in[79:72] ? 8'hf : _GEN_2298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2300 = 8'hfc == io_data_in[79:72] ? 8'hb0 : _GEN_2299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2301 = 8'hfd == io_data_in[79:72] ? 8'h54 : _GEN_2300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2302 = 8'hfe == io_data_in[79:72] ? 8'hbb : _GEN_2301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2303 = 8'hff == io_data_in[79:72] ? 8'h16 : _GEN_2302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2305 = 8'h1 == io_data_in[71:64] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2306 = 8'h2 == io_data_in[71:64] ? 8'h77 : _GEN_2305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2307 = 8'h3 == io_data_in[71:64] ? 8'h7b : _GEN_2306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2308 = 8'h4 == io_data_in[71:64] ? 8'hf2 : _GEN_2307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2309 = 8'h5 == io_data_in[71:64] ? 8'h6b : _GEN_2308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2310 = 8'h6 == io_data_in[71:64] ? 8'h6f : _GEN_2309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2311 = 8'h7 == io_data_in[71:64] ? 8'hc5 : _GEN_2310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2312 = 8'h8 == io_data_in[71:64] ? 8'h30 : _GEN_2311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2313 = 8'h9 == io_data_in[71:64] ? 8'h1 : _GEN_2312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2314 = 8'ha == io_data_in[71:64] ? 8'h67 : _GEN_2313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2315 = 8'hb == io_data_in[71:64] ? 8'h2b : _GEN_2314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2316 = 8'hc == io_data_in[71:64] ? 8'hfe : _GEN_2315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2317 = 8'hd == io_data_in[71:64] ? 8'hd7 : _GEN_2316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2318 = 8'he == io_data_in[71:64] ? 8'hab : _GEN_2317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2319 = 8'hf == io_data_in[71:64] ? 8'h76 : _GEN_2318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2320 = 8'h10 == io_data_in[71:64] ? 8'hca : _GEN_2319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2321 = 8'h11 == io_data_in[71:64] ? 8'h82 : _GEN_2320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2322 = 8'h12 == io_data_in[71:64] ? 8'hc9 : _GEN_2321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2323 = 8'h13 == io_data_in[71:64] ? 8'h7d : _GEN_2322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2324 = 8'h14 == io_data_in[71:64] ? 8'hfa : _GEN_2323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2325 = 8'h15 == io_data_in[71:64] ? 8'h59 : _GEN_2324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2326 = 8'h16 == io_data_in[71:64] ? 8'h47 : _GEN_2325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2327 = 8'h17 == io_data_in[71:64] ? 8'hf0 : _GEN_2326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2328 = 8'h18 == io_data_in[71:64] ? 8'had : _GEN_2327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2329 = 8'h19 == io_data_in[71:64] ? 8'hd4 : _GEN_2328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2330 = 8'h1a == io_data_in[71:64] ? 8'ha2 : _GEN_2329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2331 = 8'h1b == io_data_in[71:64] ? 8'haf : _GEN_2330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2332 = 8'h1c == io_data_in[71:64] ? 8'h9c : _GEN_2331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2333 = 8'h1d == io_data_in[71:64] ? 8'ha4 : _GEN_2332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2334 = 8'h1e == io_data_in[71:64] ? 8'h72 : _GEN_2333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2335 = 8'h1f == io_data_in[71:64] ? 8'hc0 : _GEN_2334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2336 = 8'h20 == io_data_in[71:64] ? 8'hb7 : _GEN_2335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2337 = 8'h21 == io_data_in[71:64] ? 8'hfd : _GEN_2336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2338 = 8'h22 == io_data_in[71:64] ? 8'h93 : _GEN_2337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2339 = 8'h23 == io_data_in[71:64] ? 8'h26 : _GEN_2338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2340 = 8'h24 == io_data_in[71:64] ? 8'h36 : _GEN_2339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2341 = 8'h25 == io_data_in[71:64] ? 8'h3f : _GEN_2340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2342 = 8'h26 == io_data_in[71:64] ? 8'hf7 : _GEN_2341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2343 = 8'h27 == io_data_in[71:64] ? 8'hcc : _GEN_2342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2344 = 8'h28 == io_data_in[71:64] ? 8'h34 : _GEN_2343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2345 = 8'h29 == io_data_in[71:64] ? 8'ha5 : _GEN_2344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2346 = 8'h2a == io_data_in[71:64] ? 8'he5 : _GEN_2345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2347 = 8'h2b == io_data_in[71:64] ? 8'hf1 : _GEN_2346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2348 = 8'h2c == io_data_in[71:64] ? 8'h71 : _GEN_2347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2349 = 8'h2d == io_data_in[71:64] ? 8'hd8 : _GEN_2348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2350 = 8'h2e == io_data_in[71:64] ? 8'h31 : _GEN_2349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2351 = 8'h2f == io_data_in[71:64] ? 8'h15 : _GEN_2350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2352 = 8'h30 == io_data_in[71:64] ? 8'h4 : _GEN_2351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2353 = 8'h31 == io_data_in[71:64] ? 8'hc7 : _GEN_2352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2354 = 8'h32 == io_data_in[71:64] ? 8'h23 : _GEN_2353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2355 = 8'h33 == io_data_in[71:64] ? 8'hc3 : _GEN_2354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2356 = 8'h34 == io_data_in[71:64] ? 8'h18 : _GEN_2355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2357 = 8'h35 == io_data_in[71:64] ? 8'h96 : _GEN_2356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2358 = 8'h36 == io_data_in[71:64] ? 8'h5 : _GEN_2357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2359 = 8'h37 == io_data_in[71:64] ? 8'h9a : _GEN_2358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2360 = 8'h38 == io_data_in[71:64] ? 8'h7 : _GEN_2359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2361 = 8'h39 == io_data_in[71:64] ? 8'h12 : _GEN_2360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2362 = 8'h3a == io_data_in[71:64] ? 8'h80 : _GEN_2361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2363 = 8'h3b == io_data_in[71:64] ? 8'he2 : _GEN_2362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2364 = 8'h3c == io_data_in[71:64] ? 8'heb : _GEN_2363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2365 = 8'h3d == io_data_in[71:64] ? 8'h27 : _GEN_2364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2366 = 8'h3e == io_data_in[71:64] ? 8'hb2 : _GEN_2365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2367 = 8'h3f == io_data_in[71:64] ? 8'h75 : _GEN_2366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2368 = 8'h40 == io_data_in[71:64] ? 8'h9 : _GEN_2367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2369 = 8'h41 == io_data_in[71:64] ? 8'h83 : _GEN_2368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2370 = 8'h42 == io_data_in[71:64] ? 8'h2c : _GEN_2369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2371 = 8'h43 == io_data_in[71:64] ? 8'h1a : _GEN_2370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2372 = 8'h44 == io_data_in[71:64] ? 8'h1b : _GEN_2371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2373 = 8'h45 == io_data_in[71:64] ? 8'h6e : _GEN_2372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2374 = 8'h46 == io_data_in[71:64] ? 8'h5a : _GEN_2373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2375 = 8'h47 == io_data_in[71:64] ? 8'ha0 : _GEN_2374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2376 = 8'h48 == io_data_in[71:64] ? 8'h52 : _GEN_2375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2377 = 8'h49 == io_data_in[71:64] ? 8'h3b : _GEN_2376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2378 = 8'h4a == io_data_in[71:64] ? 8'hd6 : _GEN_2377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2379 = 8'h4b == io_data_in[71:64] ? 8'hb3 : _GEN_2378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2380 = 8'h4c == io_data_in[71:64] ? 8'h29 : _GEN_2379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2381 = 8'h4d == io_data_in[71:64] ? 8'he3 : _GEN_2380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2382 = 8'h4e == io_data_in[71:64] ? 8'h2f : _GEN_2381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2383 = 8'h4f == io_data_in[71:64] ? 8'h84 : _GEN_2382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2384 = 8'h50 == io_data_in[71:64] ? 8'h53 : _GEN_2383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2385 = 8'h51 == io_data_in[71:64] ? 8'hd1 : _GEN_2384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2386 = 8'h52 == io_data_in[71:64] ? 8'h0 : _GEN_2385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2387 = 8'h53 == io_data_in[71:64] ? 8'hed : _GEN_2386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2388 = 8'h54 == io_data_in[71:64] ? 8'h20 : _GEN_2387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2389 = 8'h55 == io_data_in[71:64] ? 8'hfc : _GEN_2388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2390 = 8'h56 == io_data_in[71:64] ? 8'hb1 : _GEN_2389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2391 = 8'h57 == io_data_in[71:64] ? 8'h5b : _GEN_2390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2392 = 8'h58 == io_data_in[71:64] ? 8'h6a : _GEN_2391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2393 = 8'h59 == io_data_in[71:64] ? 8'hcb : _GEN_2392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2394 = 8'h5a == io_data_in[71:64] ? 8'hbe : _GEN_2393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2395 = 8'h5b == io_data_in[71:64] ? 8'h39 : _GEN_2394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2396 = 8'h5c == io_data_in[71:64] ? 8'h4a : _GEN_2395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2397 = 8'h5d == io_data_in[71:64] ? 8'h4c : _GEN_2396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2398 = 8'h5e == io_data_in[71:64] ? 8'h58 : _GEN_2397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2399 = 8'h5f == io_data_in[71:64] ? 8'hcf : _GEN_2398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2400 = 8'h60 == io_data_in[71:64] ? 8'hd0 : _GEN_2399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2401 = 8'h61 == io_data_in[71:64] ? 8'hef : _GEN_2400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2402 = 8'h62 == io_data_in[71:64] ? 8'haa : _GEN_2401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2403 = 8'h63 == io_data_in[71:64] ? 8'hfb : _GEN_2402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2404 = 8'h64 == io_data_in[71:64] ? 8'h43 : _GEN_2403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2405 = 8'h65 == io_data_in[71:64] ? 8'h4d : _GEN_2404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2406 = 8'h66 == io_data_in[71:64] ? 8'h33 : _GEN_2405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2407 = 8'h67 == io_data_in[71:64] ? 8'h85 : _GEN_2406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2408 = 8'h68 == io_data_in[71:64] ? 8'h45 : _GEN_2407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2409 = 8'h69 == io_data_in[71:64] ? 8'hf9 : _GEN_2408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2410 = 8'h6a == io_data_in[71:64] ? 8'h2 : _GEN_2409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2411 = 8'h6b == io_data_in[71:64] ? 8'h7f : _GEN_2410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2412 = 8'h6c == io_data_in[71:64] ? 8'h50 : _GEN_2411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2413 = 8'h6d == io_data_in[71:64] ? 8'h3c : _GEN_2412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2414 = 8'h6e == io_data_in[71:64] ? 8'h9f : _GEN_2413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2415 = 8'h6f == io_data_in[71:64] ? 8'ha8 : _GEN_2414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2416 = 8'h70 == io_data_in[71:64] ? 8'h51 : _GEN_2415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2417 = 8'h71 == io_data_in[71:64] ? 8'ha3 : _GEN_2416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2418 = 8'h72 == io_data_in[71:64] ? 8'h40 : _GEN_2417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2419 = 8'h73 == io_data_in[71:64] ? 8'h8f : _GEN_2418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2420 = 8'h74 == io_data_in[71:64] ? 8'h92 : _GEN_2419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2421 = 8'h75 == io_data_in[71:64] ? 8'h9d : _GEN_2420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2422 = 8'h76 == io_data_in[71:64] ? 8'h38 : _GEN_2421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2423 = 8'h77 == io_data_in[71:64] ? 8'hf5 : _GEN_2422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2424 = 8'h78 == io_data_in[71:64] ? 8'hbc : _GEN_2423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2425 = 8'h79 == io_data_in[71:64] ? 8'hb6 : _GEN_2424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2426 = 8'h7a == io_data_in[71:64] ? 8'hda : _GEN_2425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2427 = 8'h7b == io_data_in[71:64] ? 8'h21 : _GEN_2426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2428 = 8'h7c == io_data_in[71:64] ? 8'h10 : _GEN_2427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2429 = 8'h7d == io_data_in[71:64] ? 8'hff : _GEN_2428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2430 = 8'h7e == io_data_in[71:64] ? 8'hf3 : _GEN_2429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2431 = 8'h7f == io_data_in[71:64] ? 8'hd2 : _GEN_2430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2432 = 8'h80 == io_data_in[71:64] ? 8'hcd : _GEN_2431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2433 = 8'h81 == io_data_in[71:64] ? 8'hc : _GEN_2432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2434 = 8'h82 == io_data_in[71:64] ? 8'h13 : _GEN_2433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2435 = 8'h83 == io_data_in[71:64] ? 8'hec : _GEN_2434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2436 = 8'h84 == io_data_in[71:64] ? 8'h5f : _GEN_2435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2437 = 8'h85 == io_data_in[71:64] ? 8'h97 : _GEN_2436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2438 = 8'h86 == io_data_in[71:64] ? 8'h44 : _GEN_2437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2439 = 8'h87 == io_data_in[71:64] ? 8'h17 : _GEN_2438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2440 = 8'h88 == io_data_in[71:64] ? 8'hc4 : _GEN_2439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2441 = 8'h89 == io_data_in[71:64] ? 8'ha7 : _GEN_2440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2442 = 8'h8a == io_data_in[71:64] ? 8'h7e : _GEN_2441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2443 = 8'h8b == io_data_in[71:64] ? 8'h3d : _GEN_2442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2444 = 8'h8c == io_data_in[71:64] ? 8'h64 : _GEN_2443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2445 = 8'h8d == io_data_in[71:64] ? 8'h5d : _GEN_2444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2446 = 8'h8e == io_data_in[71:64] ? 8'h19 : _GEN_2445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2447 = 8'h8f == io_data_in[71:64] ? 8'h73 : _GEN_2446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2448 = 8'h90 == io_data_in[71:64] ? 8'h60 : _GEN_2447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2449 = 8'h91 == io_data_in[71:64] ? 8'h81 : _GEN_2448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2450 = 8'h92 == io_data_in[71:64] ? 8'h4f : _GEN_2449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2451 = 8'h93 == io_data_in[71:64] ? 8'hdc : _GEN_2450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2452 = 8'h94 == io_data_in[71:64] ? 8'h22 : _GEN_2451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2453 = 8'h95 == io_data_in[71:64] ? 8'h2a : _GEN_2452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2454 = 8'h96 == io_data_in[71:64] ? 8'h90 : _GEN_2453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2455 = 8'h97 == io_data_in[71:64] ? 8'h88 : _GEN_2454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2456 = 8'h98 == io_data_in[71:64] ? 8'h46 : _GEN_2455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2457 = 8'h99 == io_data_in[71:64] ? 8'hee : _GEN_2456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2458 = 8'h9a == io_data_in[71:64] ? 8'hb8 : _GEN_2457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2459 = 8'h9b == io_data_in[71:64] ? 8'h14 : _GEN_2458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2460 = 8'h9c == io_data_in[71:64] ? 8'hde : _GEN_2459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2461 = 8'h9d == io_data_in[71:64] ? 8'h5e : _GEN_2460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2462 = 8'h9e == io_data_in[71:64] ? 8'hb : _GEN_2461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2463 = 8'h9f == io_data_in[71:64] ? 8'hdb : _GEN_2462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2464 = 8'ha0 == io_data_in[71:64] ? 8'he0 : _GEN_2463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2465 = 8'ha1 == io_data_in[71:64] ? 8'h32 : _GEN_2464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2466 = 8'ha2 == io_data_in[71:64] ? 8'h3a : _GEN_2465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2467 = 8'ha3 == io_data_in[71:64] ? 8'ha : _GEN_2466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2468 = 8'ha4 == io_data_in[71:64] ? 8'h49 : _GEN_2467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2469 = 8'ha5 == io_data_in[71:64] ? 8'h6 : _GEN_2468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2470 = 8'ha6 == io_data_in[71:64] ? 8'h24 : _GEN_2469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2471 = 8'ha7 == io_data_in[71:64] ? 8'h5c : _GEN_2470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2472 = 8'ha8 == io_data_in[71:64] ? 8'hc2 : _GEN_2471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2473 = 8'ha9 == io_data_in[71:64] ? 8'hd3 : _GEN_2472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2474 = 8'haa == io_data_in[71:64] ? 8'hac : _GEN_2473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2475 = 8'hab == io_data_in[71:64] ? 8'h62 : _GEN_2474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2476 = 8'hac == io_data_in[71:64] ? 8'h91 : _GEN_2475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2477 = 8'had == io_data_in[71:64] ? 8'h95 : _GEN_2476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2478 = 8'hae == io_data_in[71:64] ? 8'he4 : _GEN_2477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2479 = 8'haf == io_data_in[71:64] ? 8'h79 : _GEN_2478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2480 = 8'hb0 == io_data_in[71:64] ? 8'he7 : _GEN_2479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2481 = 8'hb1 == io_data_in[71:64] ? 8'hc8 : _GEN_2480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2482 = 8'hb2 == io_data_in[71:64] ? 8'h37 : _GEN_2481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2483 = 8'hb3 == io_data_in[71:64] ? 8'h6d : _GEN_2482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2484 = 8'hb4 == io_data_in[71:64] ? 8'h8d : _GEN_2483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2485 = 8'hb5 == io_data_in[71:64] ? 8'hd5 : _GEN_2484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2486 = 8'hb6 == io_data_in[71:64] ? 8'h4e : _GEN_2485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2487 = 8'hb7 == io_data_in[71:64] ? 8'ha9 : _GEN_2486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2488 = 8'hb8 == io_data_in[71:64] ? 8'h6c : _GEN_2487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2489 = 8'hb9 == io_data_in[71:64] ? 8'h56 : _GEN_2488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2490 = 8'hba == io_data_in[71:64] ? 8'hf4 : _GEN_2489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2491 = 8'hbb == io_data_in[71:64] ? 8'hea : _GEN_2490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2492 = 8'hbc == io_data_in[71:64] ? 8'h65 : _GEN_2491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2493 = 8'hbd == io_data_in[71:64] ? 8'h7a : _GEN_2492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2494 = 8'hbe == io_data_in[71:64] ? 8'hae : _GEN_2493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2495 = 8'hbf == io_data_in[71:64] ? 8'h8 : _GEN_2494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2496 = 8'hc0 == io_data_in[71:64] ? 8'hba : _GEN_2495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2497 = 8'hc1 == io_data_in[71:64] ? 8'h78 : _GEN_2496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2498 = 8'hc2 == io_data_in[71:64] ? 8'h25 : _GEN_2497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2499 = 8'hc3 == io_data_in[71:64] ? 8'h2e : _GEN_2498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2500 = 8'hc4 == io_data_in[71:64] ? 8'h1c : _GEN_2499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2501 = 8'hc5 == io_data_in[71:64] ? 8'ha6 : _GEN_2500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2502 = 8'hc6 == io_data_in[71:64] ? 8'hb4 : _GEN_2501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2503 = 8'hc7 == io_data_in[71:64] ? 8'hc6 : _GEN_2502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2504 = 8'hc8 == io_data_in[71:64] ? 8'he8 : _GEN_2503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2505 = 8'hc9 == io_data_in[71:64] ? 8'hdd : _GEN_2504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2506 = 8'hca == io_data_in[71:64] ? 8'h74 : _GEN_2505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2507 = 8'hcb == io_data_in[71:64] ? 8'h1f : _GEN_2506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2508 = 8'hcc == io_data_in[71:64] ? 8'h4b : _GEN_2507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2509 = 8'hcd == io_data_in[71:64] ? 8'hbd : _GEN_2508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2510 = 8'hce == io_data_in[71:64] ? 8'h8b : _GEN_2509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2511 = 8'hcf == io_data_in[71:64] ? 8'h8a : _GEN_2510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2512 = 8'hd0 == io_data_in[71:64] ? 8'h70 : _GEN_2511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2513 = 8'hd1 == io_data_in[71:64] ? 8'h3e : _GEN_2512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2514 = 8'hd2 == io_data_in[71:64] ? 8'hb5 : _GEN_2513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2515 = 8'hd3 == io_data_in[71:64] ? 8'h66 : _GEN_2514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2516 = 8'hd4 == io_data_in[71:64] ? 8'h48 : _GEN_2515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2517 = 8'hd5 == io_data_in[71:64] ? 8'h3 : _GEN_2516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2518 = 8'hd6 == io_data_in[71:64] ? 8'hf6 : _GEN_2517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2519 = 8'hd7 == io_data_in[71:64] ? 8'he : _GEN_2518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2520 = 8'hd8 == io_data_in[71:64] ? 8'h61 : _GEN_2519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2521 = 8'hd9 == io_data_in[71:64] ? 8'h35 : _GEN_2520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2522 = 8'hda == io_data_in[71:64] ? 8'h57 : _GEN_2521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2523 = 8'hdb == io_data_in[71:64] ? 8'hb9 : _GEN_2522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2524 = 8'hdc == io_data_in[71:64] ? 8'h86 : _GEN_2523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2525 = 8'hdd == io_data_in[71:64] ? 8'hc1 : _GEN_2524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2526 = 8'hde == io_data_in[71:64] ? 8'h1d : _GEN_2525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2527 = 8'hdf == io_data_in[71:64] ? 8'h9e : _GEN_2526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2528 = 8'he0 == io_data_in[71:64] ? 8'he1 : _GEN_2527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2529 = 8'he1 == io_data_in[71:64] ? 8'hf8 : _GEN_2528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2530 = 8'he2 == io_data_in[71:64] ? 8'h98 : _GEN_2529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2531 = 8'he3 == io_data_in[71:64] ? 8'h11 : _GEN_2530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2532 = 8'he4 == io_data_in[71:64] ? 8'h69 : _GEN_2531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2533 = 8'he5 == io_data_in[71:64] ? 8'hd9 : _GEN_2532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2534 = 8'he6 == io_data_in[71:64] ? 8'h8e : _GEN_2533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2535 = 8'he7 == io_data_in[71:64] ? 8'h94 : _GEN_2534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2536 = 8'he8 == io_data_in[71:64] ? 8'h9b : _GEN_2535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2537 = 8'he9 == io_data_in[71:64] ? 8'h1e : _GEN_2536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2538 = 8'hea == io_data_in[71:64] ? 8'h87 : _GEN_2537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2539 = 8'heb == io_data_in[71:64] ? 8'he9 : _GEN_2538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2540 = 8'hec == io_data_in[71:64] ? 8'hce : _GEN_2539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2541 = 8'hed == io_data_in[71:64] ? 8'h55 : _GEN_2540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2542 = 8'hee == io_data_in[71:64] ? 8'h28 : _GEN_2541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2543 = 8'hef == io_data_in[71:64] ? 8'hdf : _GEN_2542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2544 = 8'hf0 == io_data_in[71:64] ? 8'h8c : _GEN_2543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2545 = 8'hf1 == io_data_in[71:64] ? 8'ha1 : _GEN_2544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2546 = 8'hf2 == io_data_in[71:64] ? 8'h89 : _GEN_2545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2547 = 8'hf3 == io_data_in[71:64] ? 8'hd : _GEN_2546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2548 = 8'hf4 == io_data_in[71:64] ? 8'hbf : _GEN_2547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2549 = 8'hf5 == io_data_in[71:64] ? 8'he6 : _GEN_2548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2550 = 8'hf6 == io_data_in[71:64] ? 8'h42 : _GEN_2549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2551 = 8'hf7 == io_data_in[71:64] ? 8'h68 : _GEN_2550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2552 = 8'hf8 == io_data_in[71:64] ? 8'h41 : _GEN_2551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2553 = 8'hf9 == io_data_in[71:64] ? 8'h99 : _GEN_2552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2554 = 8'hfa == io_data_in[71:64] ? 8'h2d : _GEN_2553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2555 = 8'hfb == io_data_in[71:64] ? 8'hf : _GEN_2554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2556 = 8'hfc == io_data_in[71:64] ? 8'hb0 : _GEN_2555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2557 = 8'hfd == io_data_in[71:64] ? 8'h54 : _GEN_2556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2558 = 8'hfe == io_data_in[71:64] ? 8'hbb : _GEN_2557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2559 = 8'hff == io_data_in[71:64] ? 8'h16 : _GEN_2558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2561 = 8'h1 == io_data_in[95:88] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2562 = 8'h2 == io_data_in[95:88] ? 8'h77 : _GEN_2561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2563 = 8'h3 == io_data_in[95:88] ? 8'h7b : _GEN_2562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2564 = 8'h4 == io_data_in[95:88] ? 8'hf2 : _GEN_2563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2565 = 8'h5 == io_data_in[95:88] ? 8'h6b : _GEN_2564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2566 = 8'h6 == io_data_in[95:88] ? 8'h6f : _GEN_2565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2567 = 8'h7 == io_data_in[95:88] ? 8'hc5 : _GEN_2566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2568 = 8'h8 == io_data_in[95:88] ? 8'h30 : _GEN_2567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2569 = 8'h9 == io_data_in[95:88] ? 8'h1 : _GEN_2568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2570 = 8'ha == io_data_in[95:88] ? 8'h67 : _GEN_2569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2571 = 8'hb == io_data_in[95:88] ? 8'h2b : _GEN_2570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2572 = 8'hc == io_data_in[95:88] ? 8'hfe : _GEN_2571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2573 = 8'hd == io_data_in[95:88] ? 8'hd7 : _GEN_2572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2574 = 8'he == io_data_in[95:88] ? 8'hab : _GEN_2573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2575 = 8'hf == io_data_in[95:88] ? 8'h76 : _GEN_2574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2576 = 8'h10 == io_data_in[95:88] ? 8'hca : _GEN_2575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2577 = 8'h11 == io_data_in[95:88] ? 8'h82 : _GEN_2576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2578 = 8'h12 == io_data_in[95:88] ? 8'hc9 : _GEN_2577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2579 = 8'h13 == io_data_in[95:88] ? 8'h7d : _GEN_2578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2580 = 8'h14 == io_data_in[95:88] ? 8'hfa : _GEN_2579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2581 = 8'h15 == io_data_in[95:88] ? 8'h59 : _GEN_2580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2582 = 8'h16 == io_data_in[95:88] ? 8'h47 : _GEN_2581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2583 = 8'h17 == io_data_in[95:88] ? 8'hf0 : _GEN_2582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2584 = 8'h18 == io_data_in[95:88] ? 8'had : _GEN_2583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2585 = 8'h19 == io_data_in[95:88] ? 8'hd4 : _GEN_2584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2586 = 8'h1a == io_data_in[95:88] ? 8'ha2 : _GEN_2585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2587 = 8'h1b == io_data_in[95:88] ? 8'haf : _GEN_2586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2588 = 8'h1c == io_data_in[95:88] ? 8'h9c : _GEN_2587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2589 = 8'h1d == io_data_in[95:88] ? 8'ha4 : _GEN_2588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2590 = 8'h1e == io_data_in[95:88] ? 8'h72 : _GEN_2589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2591 = 8'h1f == io_data_in[95:88] ? 8'hc0 : _GEN_2590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2592 = 8'h20 == io_data_in[95:88] ? 8'hb7 : _GEN_2591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2593 = 8'h21 == io_data_in[95:88] ? 8'hfd : _GEN_2592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2594 = 8'h22 == io_data_in[95:88] ? 8'h93 : _GEN_2593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2595 = 8'h23 == io_data_in[95:88] ? 8'h26 : _GEN_2594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2596 = 8'h24 == io_data_in[95:88] ? 8'h36 : _GEN_2595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2597 = 8'h25 == io_data_in[95:88] ? 8'h3f : _GEN_2596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2598 = 8'h26 == io_data_in[95:88] ? 8'hf7 : _GEN_2597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2599 = 8'h27 == io_data_in[95:88] ? 8'hcc : _GEN_2598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2600 = 8'h28 == io_data_in[95:88] ? 8'h34 : _GEN_2599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2601 = 8'h29 == io_data_in[95:88] ? 8'ha5 : _GEN_2600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2602 = 8'h2a == io_data_in[95:88] ? 8'he5 : _GEN_2601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2603 = 8'h2b == io_data_in[95:88] ? 8'hf1 : _GEN_2602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2604 = 8'h2c == io_data_in[95:88] ? 8'h71 : _GEN_2603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2605 = 8'h2d == io_data_in[95:88] ? 8'hd8 : _GEN_2604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2606 = 8'h2e == io_data_in[95:88] ? 8'h31 : _GEN_2605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2607 = 8'h2f == io_data_in[95:88] ? 8'h15 : _GEN_2606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2608 = 8'h30 == io_data_in[95:88] ? 8'h4 : _GEN_2607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2609 = 8'h31 == io_data_in[95:88] ? 8'hc7 : _GEN_2608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2610 = 8'h32 == io_data_in[95:88] ? 8'h23 : _GEN_2609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2611 = 8'h33 == io_data_in[95:88] ? 8'hc3 : _GEN_2610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2612 = 8'h34 == io_data_in[95:88] ? 8'h18 : _GEN_2611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2613 = 8'h35 == io_data_in[95:88] ? 8'h96 : _GEN_2612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2614 = 8'h36 == io_data_in[95:88] ? 8'h5 : _GEN_2613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2615 = 8'h37 == io_data_in[95:88] ? 8'h9a : _GEN_2614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2616 = 8'h38 == io_data_in[95:88] ? 8'h7 : _GEN_2615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2617 = 8'h39 == io_data_in[95:88] ? 8'h12 : _GEN_2616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2618 = 8'h3a == io_data_in[95:88] ? 8'h80 : _GEN_2617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2619 = 8'h3b == io_data_in[95:88] ? 8'he2 : _GEN_2618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2620 = 8'h3c == io_data_in[95:88] ? 8'heb : _GEN_2619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2621 = 8'h3d == io_data_in[95:88] ? 8'h27 : _GEN_2620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2622 = 8'h3e == io_data_in[95:88] ? 8'hb2 : _GEN_2621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2623 = 8'h3f == io_data_in[95:88] ? 8'h75 : _GEN_2622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2624 = 8'h40 == io_data_in[95:88] ? 8'h9 : _GEN_2623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2625 = 8'h41 == io_data_in[95:88] ? 8'h83 : _GEN_2624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2626 = 8'h42 == io_data_in[95:88] ? 8'h2c : _GEN_2625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2627 = 8'h43 == io_data_in[95:88] ? 8'h1a : _GEN_2626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2628 = 8'h44 == io_data_in[95:88] ? 8'h1b : _GEN_2627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2629 = 8'h45 == io_data_in[95:88] ? 8'h6e : _GEN_2628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2630 = 8'h46 == io_data_in[95:88] ? 8'h5a : _GEN_2629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2631 = 8'h47 == io_data_in[95:88] ? 8'ha0 : _GEN_2630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2632 = 8'h48 == io_data_in[95:88] ? 8'h52 : _GEN_2631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2633 = 8'h49 == io_data_in[95:88] ? 8'h3b : _GEN_2632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2634 = 8'h4a == io_data_in[95:88] ? 8'hd6 : _GEN_2633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2635 = 8'h4b == io_data_in[95:88] ? 8'hb3 : _GEN_2634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2636 = 8'h4c == io_data_in[95:88] ? 8'h29 : _GEN_2635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2637 = 8'h4d == io_data_in[95:88] ? 8'he3 : _GEN_2636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2638 = 8'h4e == io_data_in[95:88] ? 8'h2f : _GEN_2637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2639 = 8'h4f == io_data_in[95:88] ? 8'h84 : _GEN_2638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2640 = 8'h50 == io_data_in[95:88] ? 8'h53 : _GEN_2639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2641 = 8'h51 == io_data_in[95:88] ? 8'hd1 : _GEN_2640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2642 = 8'h52 == io_data_in[95:88] ? 8'h0 : _GEN_2641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2643 = 8'h53 == io_data_in[95:88] ? 8'hed : _GEN_2642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2644 = 8'h54 == io_data_in[95:88] ? 8'h20 : _GEN_2643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2645 = 8'h55 == io_data_in[95:88] ? 8'hfc : _GEN_2644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2646 = 8'h56 == io_data_in[95:88] ? 8'hb1 : _GEN_2645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2647 = 8'h57 == io_data_in[95:88] ? 8'h5b : _GEN_2646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2648 = 8'h58 == io_data_in[95:88] ? 8'h6a : _GEN_2647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2649 = 8'h59 == io_data_in[95:88] ? 8'hcb : _GEN_2648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2650 = 8'h5a == io_data_in[95:88] ? 8'hbe : _GEN_2649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2651 = 8'h5b == io_data_in[95:88] ? 8'h39 : _GEN_2650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2652 = 8'h5c == io_data_in[95:88] ? 8'h4a : _GEN_2651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2653 = 8'h5d == io_data_in[95:88] ? 8'h4c : _GEN_2652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2654 = 8'h5e == io_data_in[95:88] ? 8'h58 : _GEN_2653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2655 = 8'h5f == io_data_in[95:88] ? 8'hcf : _GEN_2654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2656 = 8'h60 == io_data_in[95:88] ? 8'hd0 : _GEN_2655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2657 = 8'h61 == io_data_in[95:88] ? 8'hef : _GEN_2656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2658 = 8'h62 == io_data_in[95:88] ? 8'haa : _GEN_2657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2659 = 8'h63 == io_data_in[95:88] ? 8'hfb : _GEN_2658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2660 = 8'h64 == io_data_in[95:88] ? 8'h43 : _GEN_2659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2661 = 8'h65 == io_data_in[95:88] ? 8'h4d : _GEN_2660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2662 = 8'h66 == io_data_in[95:88] ? 8'h33 : _GEN_2661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2663 = 8'h67 == io_data_in[95:88] ? 8'h85 : _GEN_2662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2664 = 8'h68 == io_data_in[95:88] ? 8'h45 : _GEN_2663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2665 = 8'h69 == io_data_in[95:88] ? 8'hf9 : _GEN_2664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2666 = 8'h6a == io_data_in[95:88] ? 8'h2 : _GEN_2665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2667 = 8'h6b == io_data_in[95:88] ? 8'h7f : _GEN_2666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2668 = 8'h6c == io_data_in[95:88] ? 8'h50 : _GEN_2667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2669 = 8'h6d == io_data_in[95:88] ? 8'h3c : _GEN_2668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2670 = 8'h6e == io_data_in[95:88] ? 8'h9f : _GEN_2669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2671 = 8'h6f == io_data_in[95:88] ? 8'ha8 : _GEN_2670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2672 = 8'h70 == io_data_in[95:88] ? 8'h51 : _GEN_2671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2673 = 8'h71 == io_data_in[95:88] ? 8'ha3 : _GEN_2672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2674 = 8'h72 == io_data_in[95:88] ? 8'h40 : _GEN_2673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2675 = 8'h73 == io_data_in[95:88] ? 8'h8f : _GEN_2674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2676 = 8'h74 == io_data_in[95:88] ? 8'h92 : _GEN_2675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2677 = 8'h75 == io_data_in[95:88] ? 8'h9d : _GEN_2676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2678 = 8'h76 == io_data_in[95:88] ? 8'h38 : _GEN_2677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2679 = 8'h77 == io_data_in[95:88] ? 8'hf5 : _GEN_2678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2680 = 8'h78 == io_data_in[95:88] ? 8'hbc : _GEN_2679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2681 = 8'h79 == io_data_in[95:88] ? 8'hb6 : _GEN_2680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2682 = 8'h7a == io_data_in[95:88] ? 8'hda : _GEN_2681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2683 = 8'h7b == io_data_in[95:88] ? 8'h21 : _GEN_2682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2684 = 8'h7c == io_data_in[95:88] ? 8'h10 : _GEN_2683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2685 = 8'h7d == io_data_in[95:88] ? 8'hff : _GEN_2684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2686 = 8'h7e == io_data_in[95:88] ? 8'hf3 : _GEN_2685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2687 = 8'h7f == io_data_in[95:88] ? 8'hd2 : _GEN_2686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2688 = 8'h80 == io_data_in[95:88] ? 8'hcd : _GEN_2687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2689 = 8'h81 == io_data_in[95:88] ? 8'hc : _GEN_2688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2690 = 8'h82 == io_data_in[95:88] ? 8'h13 : _GEN_2689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2691 = 8'h83 == io_data_in[95:88] ? 8'hec : _GEN_2690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2692 = 8'h84 == io_data_in[95:88] ? 8'h5f : _GEN_2691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2693 = 8'h85 == io_data_in[95:88] ? 8'h97 : _GEN_2692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2694 = 8'h86 == io_data_in[95:88] ? 8'h44 : _GEN_2693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2695 = 8'h87 == io_data_in[95:88] ? 8'h17 : _GEN_2694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2696 = 8'h88 == io_data_in[95:88] ? 8'hc4 : _GEN_2695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2697 = 8'h89 == io_data_in[95:88] ? 8'ha7 : _GEN_2696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2698 = 8'h8a == io_data_in[95:88] ? 8'h7e : _GEN_2697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2699 = 8'h8b == io_data_in[95:88] ? 8'h3d : _GEN_2698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2700 = 8'h8c == io_data_in[95:88] ? 8'h64 : _GEN_2699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2701 = 8'h8d == io_data_in[95:88] ? 8'h5d : _GEN_2700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2702 = 8'h8e == io_data_in[95:88] ? 8'h19 : _GEN_2701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2703 = 8'h8f == io_data_in[95:88] ? 8'h73 : _GEN_2702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2704 = 8'h90 == io_data_in[95:88] ? 8'h60 : _GEN_2703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2705 = 8'h91 == io_data_in[95:88] ? 8'h81 : _GEN_2704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2706 = 8'h92 == io_data_in[95:88] ? 8'h4f : _GEN_2705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2707 = 8'h93 == io_data_in[95:88] ? 8'hdc : _GEN_2706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2708 = 8'h94 == io_data_in[95:88] ? 8'h22 : _GEN_2707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2709 = 8'h95 == io_data_in[95:88] ? 8'h2a : _GEN_2708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2710 = 8'h96 == io_data_in[95:88] ? 8'h90 : _GEN_2709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2711 = 8'h97 == io_data_in[95:88] ? 8'h88 : _GEN_2710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2712 = 8'h98 == io_data_in[95:88] ? 8'h46 : _GEN_2711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2713 = 8'h99 == io_data_in[95:88] ? 8'hee : _GEN_2712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2714 = 8'h9a == io_data_in[95:88] ? 8'hb8 : _GEN_2713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2715 = 8'h9b == io_data_in[95:88] ? 8'h14 : _GEN_2714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2716 = 8'h9c == io_data_in[95:88] ? 8'hde : _GEN_2715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2717 = 8'h9d == io_data_in[95:88] ? 8'h5e : _GEN_2716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2718 = 8'h9e == io_data_in[95:88] ? 8'hb : _GEN_2717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2719 = 8'h9f == io_data_in[95:88] ? 8'hdb : _GEN_2718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2720 = 8'ha0 == io_data_in[95:88] ? 8'he0 : _GEN_2719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2721 = 8'ha1 == io_data_in[95:88] ? 8'h32 : _GEN_2720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2722 = 8'ha2 == io_data_in[95:88] ? 8'h3a : _GEN_2721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2723 = 8'ha3 == io_data_in[95:88] ? 8'ha : _GEN_2722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2724 = 8'ha4 == io_data_in[95:88] ? 8'h49 : _GEN_2723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2725 = 8'ha5 == io_data_in[95:88] ? 8'h6 : _GEN_2724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2726 = 8'ha6 == io_data_in[95:88] ? 8'h24 : _GEN_2725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2727 = 8'ha7 == io_data_in[95:88] ? 8'h5c : _GEN_2726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2728 = 8'ha8 == io_data_in[95:88] ? 8'hc2 : _GEN_2727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2729 = 8'ha9 == io_data_in[95:88] ? 8'hd3 : _GEN_2728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2730 = 8'haa == io_data_in[95:88] ? 8'hac : _GEN_2729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2731 = 8'hab == io_data_in[95:88] ? 8'h62 : _GEN_2730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2732 = 8'hac == io_data_in[95:88] ? 8'h91 : _GEN_2731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2733 = 8'had == io_data_in[95:88] ? 8'h95 : _GEN_2732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2734 = 8'hae == io_data_in[95:88] ? 8'he4 : _GEN_2733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2735 = 8'haf == io_data_in[95:88] ? 8'h79 : _GEN_2734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2736 = 8'hb0 == io_data_in[95:88] ? 8'he7 : _GEN_2735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2737 = 8'hb1 == io_data_in[95:88] ? 8'hc8 : _GEN_2736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2738 = 8'hb2 == io_data_in[95:88] ? 8'h37 : _GEN_2737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2739 = 8'hb3 == io_data_in[95:88] ? 8'h6d : _GEN_2738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2740 = 8'hb4 == io_data_in[95:88] ? 8'h8d : _GEN_2739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2741 = 8'hb5 == io_data_in[95:88] ? 8'hd5 : _GEN_2740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2742 = 8'hb6 == io_data_in[95:88] ? 8'h4e : _GEN_2741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2743 = 8'hb7 == io_data_in[95:88] ? 8'ha9 : _GEN_2742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2744 = 8'hb8 == io_data_in[95:88] ? 8'h6c : _GEN_2743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2745 = 8'hb9 == io_data_in[95:88] ? 8'h56 : _GEN_2744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2746 = 8'hba == io_data_in[95:88] ? 8'hf4 : _GEN_2745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2747 = 8'hbb == io_data_in[95:88] ? 8'hea : _GEN_2746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2748 = 8'hbc == io_data_in[95:88] ? 8'h65 : _GEN_2747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2749 = 8'hbd == io_data_in[95:88] ? 8'h7a : _GEN_2748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2750 = 8'hbe == io_data_in[95:88] ? 8'hae : _GEN_2749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2751 = 8'hbf == io_data_in[95:88] ? 8'h8 : _GEN_2750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2752 = 8'hc0 == io_data_in[95:88] ? 8'hba : _GEN_2751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2753 = 8'hc1 == io_data_in[95:88] ? 8'h78 : _GEN_2752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2754 = 8'hc2 == io_data_in[95:88] ? 8'h25 : _GEN_2753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2755 = 8'hc3 == io_data_in[95:88] ? 8'h2e : _GEN_2754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2756 = 8'hc4 == io_data_in[95:88] ? 8'h1c : _GEN_2755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2757 = 8'hc5 == io_data_in[95:88] ? 8'ha6 : _GEN_2756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2758 = 8'hc6 == io_data_in[95:88] ? 8'hb4 : _GEN_2757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2759 = 8'hc7 == io_data_in[95:88] ? 8'hc6 : _GEN_2758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2760 = 8'hc8 == io_data_in[95:88] ? 8'he8 : _GEN_2759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2761 = 8'hc9 == io_data_in[95:88] ? 8'hdd : _GEN_2760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2762 = 8'hca == io_data_in[95:88] ? 8'h74 : _GEN_2761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2763 = 8'hcb == io_data_in[95:88] ? 8'h1f : _GEN_2762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2764 = 8'hcc == io_data_in[95:88] ? 8'h4b : _GEN_2763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2765 = 8'hcd == io_data_in[95:88] ? 8'hbd : _GEN_2764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2766 = 8'hce == io_data_in[95:88] ? 8'h8b : _GEN_2765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2767 = 8'hcf == io_data_in[95:88] ? 8'h8a : _GEN_2766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2768 = 8'hd0 == io_data_in[95:88] ? 8'h70 : _GEN_2767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2769 = 8'hd1 == io_data_in[95:88] ? 8'h3e : _GEN_2768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2770 = 8'hd2 == io_data_in[95:88] ? 8'hb5 : _GEN_2769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2771 = 8'hd3 == io_data_in[95:88] ? 8'h66 : _GEN_2770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2772 = 8'hd4 == io_data_in[95:88] ? 8'h48 : _GEN_2771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2773 = 8'hd5 == io_data_in[95:88] ? 8'h3 : _GEN_2772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2774 = 8'hd6 == io_data_in[95:88] ? 8'hf6 : _GEN_2773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2775 = 8'hd7 == io_data_in[95:88] ? 8'he : _GEN_2774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2776 = 8'hd8 == io_data_in[95:88] ? 8'h61 : _GEN_2775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2777 = 8'hd9 == io_data_in[95:88] ? 8'h35 : _GEN_2776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2778 = 8'hda == io_data_in[95:88] ? 8'h57 : _GEN_2777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2779 = 8'hdb == io_data_in[95:88] ? 8'hb9 : _GEN_2778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2780 = 8'hdc == io_data_in[95:88] ? 8'h86 : _GEN_2779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2781 = 8'hdd == io_data_in[95:88] ? 8'hc1 : _GEN_2780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2782 = 8'hde == io_data_in[95:88] ? 8'h1d : _GEN_2781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2783 = 8'hdf == io_data_in[95:88] ? 8'h9e : _GEN_2782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2784 = 8'he0 == io_data_in[95:88] ? 8'he1 : _GEN_2783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2785 = 8'he1 == io_data_in[95:88] ? 8'hf8 : _GEN_2784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2786 = 8'he2 == io_data_in[95:88] ? 8'h98 : _GEN_2785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2787 = 8'he3 == io_data_in[95:88] ? 8'h11 : _GEN_2786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2788 = 8'he4 == io_data_in[95:88] ? 8'h69 : _GEN_2787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2789 = 8'he5 == io_data_in[95:88] ? 8'hd9 : _GEN_2788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2790 = 8'he6 == io_data_in[95:88] ? 8'h8e : _GEN_2789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2791 = 8'he7 == io_data_in[95:88] ? 8'h94 : _GEN_2790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2792 = 8'he8 == io_data_in[95:88] ? 8'h9b : _GEN_2791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2793 = 8'he9 == io_data_in[95:88] ? 8'h1e : _GEN_2792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2794 = 8'hea == io_data_in[95:88] ? 8'h87 : _GEN_2793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2795 = 8'heb == io_data_in[95:88] ? 8'he9 : _GEN_2794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2796 = 8'hec == io_data_in[95:88] ? 8'hce : _GEN_2795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2797 = 8'hed == io_data_in[95:88] ? 8'h55 : _GEN_2796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2798 = 8'hee == io_data_in[95:88] ? 8'h28 : _GEN_2797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2799 = 8'hef == io_data_in[95:88] ? 8'hdf : _GEN_2798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2800 = 8'hf0 == io_data_in[95:88] ? 8'h8c : _GEN_2799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2801 = 8'hf1 == io_data_in[95:88] ? 8'ha1 : _GEN_2800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2802 = 8'hf2 == io_data_in[95:88] ? 8'h89 : _GEN_2801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2803 = 8'hf3 == io_data_in[95:88] ? 8'hd : _GEN_2802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2804 = 8'hf4 == io_data_in[95:88] ? 8'hbf : _GEN_2803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2805 = 8'hf5 == io_data_in[95:88] ? 8'he6 : _GEN_2804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2806 = 8'hf6 == io_data_in[95:88] ? 8'h42 : _GEN_2805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2807 = 8'hf7 == io_data_in[95:88] ? 8'h68 : _GEN_2806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2808 = 8'hf8 == io_data_in[95:88] ? 8'h41 : _GEN_2807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2809 = 8'hf9 == io_data_in[95:88] ? 8'h99 : _GEN_2808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2810 = 8'hfa == io_data_in[95:88] ? 8'h2d : _GEN_2809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2811 = 8'hfb == io_data_in[95:88] ? 8'hf : _GEN_2810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2812 = 8'hfc == io_data_in[95:88] ? 8'hb0 : _GEN_2811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2813 = 8'hfd == io_data_in[95:88] ? 8'h54 : _GEN_2812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2814 = 8'hfe == io_data_in[95:88] ? 8'hbb : _GEN_2813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2815 = 8'hff == io_data_in[95:88] ? 8'h16 : _GEN_2814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2817 = 8'h1 == io_data_in[87:80] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2818 = 8'h2 == io_data_in[87:80] ? 8'h77 : _GEN_2817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2819 = 8'h3 == io_data_in[87:80] ? 8'h7b : _GEN_2818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2820 = 8'h4 == io_data_in[87:80] ? 8'hf2 : _GEN_2819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2821 = 8'h5 == io_data_in[87:80] ? 8'h6b : _GEN_2820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2822 = 8'h6 == io_data_in[87:80] ? 8'h6f : _GEN_2821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2823 = 8'h7 == io_data_in[87:80] ? 8'hc5 : _GEN_2822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2824 = 8'h8 == io_data_in[87:80] ? 8'h30 : _GEN_2823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2825 = 8'h9 == io_data_in[87:80] ? 8'h1 : _GEN_2824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2826 = 8'ha == io_data_in[87:80] ? 8'h67 : _GEN_2825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2827 = 8'hb == io_data_in[87:80] ? 8'h2b : _GEN_2826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2828 = 8'hc == io_data_in[87:80] ? 8'hfe : _GEN_2827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2829 = 8'hd == io_data_in[87:80] ? 8'hd7 : _GEN_2828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2830 = 8'he == io_data_in[87:80] ? 8'hab : _GEN_2829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2831 = 8'hf == io_data_in[87:80] ? 8'h76 : _GEN_2830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2832 = 8'h10 == io_data_in[87:80] ? 8'hca : _GEN_2831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2833 = 8'h11 == io_data_in[87:80] ? 8'h82 : _GEN_2832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2834 = 8'h12 == io_data_in[87:80] ? 8'hc9 : _GEN_2833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2835 = 8'h13 == io_data_in[87:80] ? 8'h7d : _GEN_2834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2836 = 8'h14 == io_data_in[87:80] ? 8'hfa : _GEN_2835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2837 = 8'h15 == io_data_in[87:80] ? 8'h59 : _GEN_2836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2838 = 8'h16 == io_data_in[87:80] ? 8'h47 : _GEN_2837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2839 = 8'h17 == io_data_in[87:80] ? 8'hf0 : _GEN_2838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2840 = 8'h18 == io_data_in[87:80] ? 8'had : _GEN_2839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2841 = 8'h19 == io_data_in[87:80] ? 8'hd4 : _GEN_2840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2842 = 8'h1a == io_data_in[87:80] ? 8'ha2 : _GEN_2841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2843 = 8'h1b == io_data_in[87:80] ? 8'haf : _GEN_2842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2844 = 8'h1c == io_data_in[87:80] ? 8'h9c : _GEN_2843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2845 = 8'h1d == io_data_in[87:80] ? 8'ha4 : _GEN_2844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2846 = 8'h1e == io_data_in[87:80] ? 8'h72 : _GEN_2845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2847 = 8'h1f == io_data_in[87:80] ? 8'hc0 : _GEN_2846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2848 = 8'h20 == io_data_in[87:80] ? 8'hb7 : _GEN_2847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2849 = 8'h21 == io_data_in[87:80] ? 8'hfd : _GEN_2848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2850 = 8'h22 == io_data_in[87:80] ? 8'h93 : _GEN_2849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2851 = 8'h23 == io_data_in[87:80] ? 8'h26 : _GEN_2850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2852 = 8'h24 == io_data_in[87:80] ? 8'h36 : _GEN_2851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2853 = 8'h25 == io_data_in[87:80] ? 8'h3f : _GEN_2852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2854 = 8'h26 == io_data_in[87:80] ? 8'hf7 : _GEN_2853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2855 = 8'h27 == io_data_in[87:80] ? 8'hcc : _GEN_2854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2856 = 8'h28 == io_data_in[87:80] ? 8'h34 : _GEN_2855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2857 = 8'h29 == io_data_in[87:80] ? 8'ha5 : _GEN_2856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2858 = 8'h2a == io_data_in[87:80] ? 8'he5 : _GEN_2857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2859 = 8'h2b == io_data_in[87:80] ? 8'hf1 : _GEN_2858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2860 = 8'h2c == io_data_in[87:80] ? 8'h71 : _GEN_2859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2861 = 8'h2d == io_data_in[87:80] ? 8'hd8 : _GEN_2860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2862 = 8'h2e == io_data_in[87:80] ? 8'h31 : _GEN_2861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2863 = 8'h2f == io_data_in[87:80] ? 8'h15 : _GEN_2862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2864 = 8'h30 == io_data_in[87:80] ? 8'h4 : _GEN_2863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2865 = 8'h31 == io_data_in[87:80] ? 8'hc7 : _GEN_2864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2866 = 8'h32 == io_data_in[87:80] ? 8'h23 : _GEN_2865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2867 = 8'h33 == io_data_in[87:80] ? 8'hc3 : _GEN_2866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2868 = 8'h34 == io_data_in[87:80] ? 8'h18 : _GEN_2867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2869 = 8'h35 == io_data_in[87:80] ? 8'h96 : _GEN_2868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2870 = 8'h36 == io_data_in[87:80] ? 8'h5 : _GEN_2869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2871 = 8'h37 == io_data_in[87:80] ? 8'h9a : _GEN_2870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2872 = 8'h38 == io_data_in[87:80] ? 8'h7 : _GEN_2871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2873 = 8'h39 == io_data_in[87:80] ? 8'h12 : _GEN_2872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2874 = 8'h3a == io_data_in[87:80] ? 8'h80 : _GEN_2873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2875 = 8'h3b == io_data_in[87:80] ? 8'he2 : _GEN_2874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2876 = 8'h3c == io_data_in[87:80] ? 8'heb : _GEN_2875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2877 = 8'h3d == io_data_in[87:80] ? 8'h27 : _GEN_2876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2878 = 8'h3e == io_data_in[87:80] ? 8'hb2 : _GEN_2877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2879 = 8'h3f == io_data_in[87:80] ? 8'h75 : _GEN_2878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2880 = 8'h40 == io_data_in[87:80] ? 8'h9 : _GEN_2879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2881 = 8'h41 == io_data_in[87:80] ? 8'h83 : _GEN_2880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2882 = 8'h42 == io_data_in[87:80] ? 8'h2c : _GEN_2881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2883 = 8'h43 == io_data_in[87:80] ? 8'h1a : _GEN_2882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2884 = 8'h44 == io_data_in[87:80] ? 8'h1b : _GEN_2883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2885 = 8'h45 == io_data_in[87:80] ? 8'h6e : _GEN_2884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2886 = 8'h46 == io_data_in[87:80] ? 8'h5a : _GEN_2885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2887 = 8'h47 == io_data_in[87:80] ? 8'ha0 : _GEN_2886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2888 = 8'h48 == io_data_in[87:80] ? 8'h52 : _GEN_2887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2889 = 8'h49 == io_data_in[87:80] ? 8'h3b : _GEN_2888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2890 = 8'h4a == io_data_in[87:80] ? 8'hd6 : _GEN_2889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2891 = 8'h4b == io_data_in[87:80] ? 8'hb3 : _GEN_2890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2892 = 8'h4c == io_data_in[87:80] ? 8'h29 : _GEN_2891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2893 = 8'h4d == io_data_in[87:80] ? 8'he3 : _GEN_2892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2894 = 8'h4e == io_data_in[87:80] ? 8'h2f : _GEN_2893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2895 = 8'h4f == io_data_in[87:80] ? 8'h84 : _GEN_2894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2896 = 8'h50 == io_data_in[87:80] ? 8'h53 : _GEN_2895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2897 = 8'h51 == io_data_in[87:80] ? 8'hd1 : _GEN_2896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2898 = 8'h52 == io_data_in[87:80] ? 8'h0 : _GEN_2897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2899 = 8'h53 == io_data_in[87:80] ? 8'hed : _GEN_2898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2900 = 8'h54 == io_data_in[87:80] ? 8'h20 : _GEN_2899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2901 = 8'h55 == io_data_in[87:80] ? 8'hfc : _GEN_2900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2902 = 8'h56 == io_data_in[87:80] ? 8'hb1 : _GEN_2901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2903 = 8'h57 == io_data_in[87:80] ? 8'h5b : _GEN_2902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2904 = 8'h58 == io_data_in[87:80] ? 8'h6a : _GEN_2903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2905 = 8'h59 == io_data_in[87:80] ? 8'hcb : _GEN_2904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2906 = 8'h5a == io_data_in[87:80] ? 8'hbe : _GEN_2905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2907 = 8'h5b == io_data_in[87:80] ? 8'h39 : _GEN_2906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2908 = 8'h5c == io_data_in[87:80] ? 8'h4a : _GEN_2907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2909 = 8'h5d == io_data_in[87:80] ? 8'h4c : _GEN_2908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2910 = 8'h5e == io_data_in[87:80] ? 8'h58 : _GEN_2909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2911 = 8'h5f == io_data_in[87:80] ? 8'hcf : _GEN_2910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2912 = 8'h60 == io_data_in[87:80] ? 8'hd0 : _GEN_2911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2913 = 8'h61 == io_data_in[87:80] ? 8'hef : _GEN_2912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2914 = 8'h62 == io_data_in[87:80] ? 8'haa : _GEN_2913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2915 = 8'h63 == io_data_in[87:80] ? 8'hfb : _GEN_2914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2916 = 8'h64 == io_data_in[87:80] ? 8'h43 : _GEN_2915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2917 = 8'h65 == io_data_in[87:80] ? 8'h4d : _GEN_2916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2918 = 8'h66 == io_data_in[87:80] ? 8'h33 : _GEN_2917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2919 = 8'h67 == io_data_in[87:80] ? 8'h85 : _GEN_2918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2920 = 8'h68 == io_data_in[87:80] ? 8'h45 : _GEN_2919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2921 = 8'h69 == io_data_in[87:80] ? 8'hf9 : _GEN_2920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2922 = 8'h6a == io_data_in[87:80] ? 8'h2 : _GEN_2921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2923 = 8'h6b == io_data_in[87:80] ? 8'h7f : _GEN_2922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2924 = 8'h6c == io_data_in[87:80] ? 8'h50 : _GEN_2923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2925 = 8'h6d == io_data_in[87:80] ? 8'h3c : _GEN_2924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2926 = 8'h6e == io_data_in[87:80] ? 8'h9f : _GEN_2925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2927 = 8'h6f == io_data_in[87:80] ? 8'ha8 : _GEN_2926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2928 = 8'h70 == io_data_in[87:80] ? 8'h51 : _GEN_2927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2929 = 8'h71 == io_data_in[87:80] ? 8'ha3 : _GEN_2928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2930 = 8'h72 == io_data_in[87:80] ? 8'h40 : _GEN_2929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2931 = 8'h73 == io_data_in[87:80] ? 8'h8f : _GEN_2930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2932 = 8'h74 == io_data_in[87:80] ? 8'h92 : _GEN_2931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2933 = 8'h75 == io_data_in[87:80] ? 8'h9d : _GEN_2932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2934 = 8'h76 == io_data_in[87:80] ? 8'h38 : _GEN_2933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2935 = 8'h77 == io_data_in[87:80] ? 8'hf5 : _GEN_2934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2936 = 8'h78 == io_data_in[87:80] ? 8'hbc : _GEN_2935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2937 = 8'h79 == io_data_in[87:80] ? 8'hb6 : _GEN_2936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2938 = 8'h7a == io_data_in[87:80] ? 8'hda : _GEN_2937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2939 = 8'h7b == io_data_in[87:80] ? 8'h21 : _GEN_2938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2940 = 8'h7c == io_data_in[87:80] ? 8'h10 : _GEN_2939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2941 = 8'h7d == io_data_in[87:80] ? 8'hff : _GEN_2940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2942 = 8'h7e == io_data_in[87:80] ? 8'hf3 : _GEN_2941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2943 = 8'h7f == io_data_in[87:80] ? 8'hd2 : _GEN_2942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2944 = 8'h80 == io_data_in[87:80] ? 8'hcd : _GEN_2943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2945 = 8'h81 == io_data_in[87:80] ? 8'hc : _GEN_2944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2946 = 8'h82 == io_data_in[87:80] ? 8'h13 : _GEN_2945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2947 = 8'h83 == io_data_in[87:80] ? 8'hec : _GEN_2946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2948 = 8'h84 == io_data_in[87:80] ? 8'h5f : _GEN_2947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2949 = 8'h85 == io_data_in[87:80] ? 8'h97 : _GEN_2948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2950 = 8'h86 == io_data_in[87:80] ? 8'h44 : _GEN_2949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2951 = 8'h87 == io_data_in[87:80] ? 8'h17 : _GEN_2950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2952 = 8'h88 == io_data_in[87:80] ? 8'hc4 : _GEN_2951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2953 = 8'h89 == io_data_in[87:80] ? 8'ha7 : _GEN_2952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2954 = 8'h8a == io_data_in[87:80] ? 8'h7e : _GEN_2953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2955 = 8'h8b == io_data_in[87:80] ? 8'h3d : _GEN_2954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2956 = 8'h8c == io_data_in[87:80] ? 8'h64 : _GEN_2955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2957 = 8'h8d == io_data_in[87:80] ? 8'h5d : _GEN_2956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2958 = 8'h8e == io_data_in[87:80] ? 8'h19 : _GEN_2957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2959 = 8'h8f == io_data_in[87:80] ? 8'h73 : _GEN_2958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2960 = 8'h90 == io_data_in[87:80] ? 8'h60 : _GEN_2959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2961 = 8'h91 == io_data_in[87:80] ? 8'h81 : _GEN_2960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2962 = 8'h92 == io_data_in[87:80] ? 8'h4f : _GEN_2961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2963 = 8'h93 == io_data_in[87:80] ? 8'hdc : _GEN_2962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2964 = 8'h94 == io_data_in[87:80] ? 8'h22 : _GEN_2963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2965 = 8'h95 == io_data_in[87:80] ? 8'h2a : _GEN_2964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2966 = 8'h96 == io_data_in[87:80] ? 8'h90 : _GEN_2965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2967 = 8'h97 == io_data_in[87:80] ? 8'h88 : _GEN_2966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2968 = 8'h98 == io_data_in[87:80] ? 8'h46 : _GEN_2967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2969 = 8'h99 == io_data_in[87:80] ? 8'hee : _GEN_2968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2970 = 8'h9a == io_data_in[87:80] ? 8'hb8 : _GEN_2969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2971 = 8'h9b == io_data_in[87:80] ? 8'h14 : _GEN_2970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2972 = 8'h9c == io_data_in[87:80] ? 8'hde : _GEN_2971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2973 = 8'h9d == io_data_in[87:80] ? 8'h5e : _GEN_2972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2974 = 8'h9e == io_data_in[87:80] ? 8'hb : _GEN_2973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2975 = 8'h9f == io_data_in[87:80] ? 8'hdb : _GEN_2974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2976 = 8'ha0 == io_data_in[87:80] ? 8'he0 : _GEN_2975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2977 = 8'ha1 == io_data_in[87:80] ? 8'h32 : _GEN_2976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2978 = 8'ha2 == io_data_in[87:80] ? 8'h3a : _GEN_2977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2979 = 8'ha3 == io_data_in[87:80] ? 8'ha : _GEN_2978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2980 = 8'ha4 == io_data_in[87:80] ? 8'h49 : _GEN_2979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2981 = 8'ha5 == io_data_in[87:80] ? 8'h6 : _GEN_2980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2982 = 8'ha6 == io_data_in[87:80] ? 8'h24 : _GEN_2981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2983 = 8'ha7 == io_data_in[87:80] ? 8'h5c : _GEN_2982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2984 = 8'ha8 == io_data_in[87:80] ? 8'hc2 : _GEN_2983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2985 = 8'ha9 == io_data_in[87:80] ? 8'hd3 : _GEN_2984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2986 = 8'haa == io_data_in[87:80] ? 8'hac : _GEN_2985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2987 = 8'hab == io_data_in[87:80] ? 8'h62 : _GEN_2986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2988 = 8'hac == io_data_in[87:80] ? 8'h91 : _GEN_2987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2989 = 8'had == io_data_in[87:80] ? 8'h95 : _GEN_2988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2990 = 8'hae == io_data_in[87:80] ? 8'he4 : _GEN_2989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2991 = 8'haf == io_data_in[87:80] ? 8'h79 : _GEN_2990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2992 = 8'hb0 == io_data_in[87:80] ? 8'he7 : _GEN_2991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2993 = 8'hb1 == io_data_in[87:80] ? 8'hc8 : _GEN_2992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2994 = 8'hb2 == io_data_in[87:80] ? 8'h37 : _GEN_2993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2995 = 8'hb3 == io_data_in[87:80] ? 8'h6d : _GEN_2994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2996 = 8'hb4 == io_data_in[87:80] ? 8'h8d : _GEN_2995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2997 = 8'hb5 == io_data_in[87:80] ? 8'hd5 : _GEN_2996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2998 = 8'hb6 == io_data_in[87:80] ? 8'h4e : _GEN_2997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2999 = 8'hb7 == io_data_in[87:80] ? 8'ha9 : _GEN_2998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3000 = 8'hb8 == io_data_in[87:80] ? 8'h6c : _GEN_2999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3001 = 8'hb9 == io_data_in[87:80] ? 8'h56 : _GEN_3000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3002 = 8'hba == io_data_in[87:80] ? 8'hf4 : _GEN_3001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3003 = 8'hbb == io_data_in[87:80] ? 8'hea : _GEN_3002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3004 = 8'hbc == io_data_in[87:80] ? 8'h65 : _GEN_3003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3005 = 8'hbd == io_data_in[87:80] ? 8'h7a : _GEN_3004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3006 = 8'hbe == io_data_in[87:80] ? 8'hae : _GEN_3005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3007 = 8'hbf == io_data_in[87:80] ? 8'h8 : _GEN_3006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3008 = 8'hc0 == io_data_in[87:80] ? 8'hba : _GEN_3007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3009 = 8'hc1 == io_data_in[87:80] ? 8'h78 : _GEN_3008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3010 = 8'hc2 == io_data_in[87:80] ? 8'h25 : _GEN_3009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3011 = 8'hc3 == io_data_in[87:80] ? 8'h2e : _GEN_3010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3012 = 8'hc4 == io_data_in[87:80] ? 8'h1c : _GEN_3011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3013 = 8'hc5 == io_data_in[87:80] ? 8'ha6 : _GEN_3012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3014 = 8'hc6 == io_data_in[87:80] ? 8'hb4 : _GEN_3013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3015 = 8'hc7 == io_data_in[87:80] ? 8'hc6 : _GEN_3014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3016 = 8'hc8 == io_data_in[87:80] ? 8'he8 : _GEN_3015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3017 = 8'hc9 == io_data_in[87:80] ? 8'hdd : _GEN_3016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3018 = 8'hca == io_data_in[87:80] ? 8'h74 : _GEN_3017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3019 = 8'hcb == io_data_in[87:80] ? 8'h1f : _GEN_3018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3020 = 8'hcc == io_data_in[87:80] ? 8'h4b : _GEN_3019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3021 = 8'hcd == io_data_in[87:80] ? 8'hbd : _GEN_3020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3022 = 8'hce == io_data_in[87:80] ? 8'h8b : _GEN_3021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3023 = 8'hcf == io_data_in[87:80] ? 8'h8a : _GEN_3022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3024 = 8'hd0 == io_data_in[87:80] ? 8'h70 : _GEN_3023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3025 = 8'hd1 == io_data_in[87:80] ? 8'h3e : _GEN_3024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3026 = 8'hd2 == io_data_in[87:80] ? 8'hb5 : _GEN_3025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3027 = 8'hd3 == io_data_in[87:80] ? 8'h66 : _GEN_3026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3028 = 8'hd4 == io_data_in[87:80] ? 8'h48 : _GEN_3027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3029 = 8'hd5 == io_data_in[87:80] ? 8'h3 : _GEN_3028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3030 = 8'hd6 == io_data_in[87:80] ? 8'hf6 : _GEN_3029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3031 = 8'hd7 == io_data_in[87:80] ? 8'he : _GEN_3030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3032 = 8'hd8 == io_data_in[87:80] ? 8'h61 : _GEN_3031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3033 = 8'hd9 == io_data_in[87:80] ? 8'h35 : _GEN_3032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3034 = 8'hda == io_data_in[87:80] ? 8'h57 : _GEN_3033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3035 = 8'hdb == io_data_in[87:80] ? 8'hb9 : _GEN_3034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3036 = 8'hdc == io_data_in[87:80] ? 8'h86 : _GEN_3035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3037 = 8'hdd == io_data_in[87:80] ? 8'hc1 : _GEN_3036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3038 = 8'hde == io_data_in[87:80] ? 8'h1d : _GEN_3037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3039 = 8'hdf == io_data_in[87:80] ? 8'h9e : _GEN_3038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3040 = 8'he0 == io_data_in[87:80] ? 8'he1 : _GEN_3039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3041 = 8'he1 == io_data_in[87:80] ? 8'hf8 : _GEN_3040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3042 = 8'he2 == io_data_in[87:80] ? 8'h98 : _GEN_3041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3043 = 8'he3 == io_data_in[87:80] ? 8'h11 : _GEN_3042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3044 = 8'he4 == io_data_in[87:80] ? 8'h69 : _GEN_3043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3045 = 8'he5 == io_data_in[87:80] ? 8'hd9 : _GEN_3044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3046 = 8'he6 == io_data_in[87:80] ? 8'h8e : _GEN_3045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3047 = 8'he7 == io_data_in[87:80] ? 8'h94 : _GEN_3046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3048 = 8'he8 == io_data_in[87:80] ? 8'h9b : _GEN_3047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3049 = 8'he9 == io_data_in[87:80] ? 8'h1e : _GEN_3048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3050 = 8'hea == io_data_in[87:80] ? 8'h87 : _GEN_3049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3051 = 8'heb == io_data_in[87:80] ? 8'he9 : _GEN_3050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3052 = 8'hec == io_data_in[87:80] ? 8'hce : _GEN_3051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3053 = 8'hed == io_data_in[87:80] ? 8'h55 : _GEN_3052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3054 = 8'hee == io_data_in[87:80] ? 8'h28 : _GEN_3053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3055 = 8'hef == io_data_in[87:80] ? 8'hdf : _GEN_3054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3056 = 8'hf0 == io_data_in[87:80] ? 8'h8c : _GEN_3055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3057 = 8'hf1 == io_data_in[87:80] ? 8'ha1 : _GEN_3056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3058 = 8'hf2 == io_data_in[87:80] ? 8'h89 : _GEN_3057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3059 = 8'hf3 == io_data_in[87:80] ? 8'hd : _GEN_3058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3060 = 8'hf4 == io_data_in[87:80] ? 8'hbf : _GEN_3059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3061 = 8'hf5 == io_data_in[87:80] ? 8'he6 : _GEN_3060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3062 = 8'hf6 == io_data_in[87:80] ? 8'h42 : _GEN_3061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3063 = 8'hf7 == io_data_in[87:80] ? 8'h68 : _GEN_3062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3064 = 8'hf8 == io_data_in[87:80] ? 8'h41 : _GEN_3063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3065 = 8'hf9 == io_data_in[87:80] ? 8'h99 : _GEN_3064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3066 = 8'hfa == io_data_in[87:80] ? 8'h2d : _GEN_3065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3067 = 8'hfb == io_data_in[87:80] ? 8'hf : _GEN_3066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3068 = 8'hfc == io_data_in[87:80] ? 8'hb0 : _GEN_3067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3069 = 8'hfd == io_data_in[87:80] ? 8'h54 : _GEN_3068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3070 = 8'hfe == io_data_in[87:80] ? 8'hbb : _GEN_3069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3071 = 8'hff == io_data_in[87:80] ? 8'h16 : _GEN_3070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3073 = 8'h1 == io_data_in[111:104] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3074 = 8'h2 == io_data_in[111:104] ? 8'h77 : _GEN_3073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3075 = 8'h3 == io_data_in[111:104] ? 8'h7b : _GEN_3074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3076 = 8'h4 == io_data_in[111:104] ? 8'hf2 : _GEN_3075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3077 = 8'h5 == io_data_in[111:104] ? 8'h6b : _GEN_3076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3078 = 8'h6 == io_data_in[111:104] ? 8'h6f : _GEN_3077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3079 = 8'h7 == io_data_in[111:104] ? 8'hc5 : _GEN_3078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3080 = 8'h8 == io_data_in[111:104] ? 8'h30 : _GEN_3079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3081 = 8'h9 == io_data_in[111:104] ? 8'h1 : _GEN_3080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3082 = 8'ha == io_data_in[111:104] ? 8'h67 : _GEN_3081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3083 = 8'hb == io_data_in[111:104] ? 8'h2b : _GEN_3082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3084 = 8'hc == io_data_in[111:104] ? 8'hfe : _GEN_3083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3085 = 8'hd == io_data_in[111:104] ? 8'hd7 : _GEN_3084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3086 = 8'he == io_data_in[111:104] ? 8'hab : _GEN_3085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3087 = 8'hf == io_data_in[111:104] ? 8'h76 : _GEN_3086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3088 = 8'h10 == io_data_in[111:104] ? 8'hca : _GEN_3087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3089 = 8'h11 == io_data_in[111:104] ? 8'h82 : _GEN_3088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3090 = 8'h12 == io_data_in[111:104] ? 8'hc9 : _GEN_3089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3091 = 8'h13 == io_data_in[111:104] ? 8'h7d : _GEN_3090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3092 = 8'h14 == io_data_in[111:104] ? 8'hfa : _GEN_3091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3093 = 8'h15 == io_data_in[111:104] ? 8'h59 : _GEN_3092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3094 = 8'h16 == io_data_in[111:104] ? 8'h47 : _GEN_3093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3095 = 8'h17 == io_data_in[111:104] ? 8'hf0 : _GEN_3094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3096 = 8'h18 == io_data_in[111:104] ? 8'had : _GEN_3095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3097 = 8'h19 == io_data_in[111:104] ? 8'hd4 : _GEN_3096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3098 = 8'h1a == io_data_in[111:104] ? 8'ha2 : _GEN_3097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3099 = 8'h1b == io_data_in[111:104] ? 8'haf : _GEN_3098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3100 = 8'h1c == io_data_in[111:104] ? 8'h9c : _GEN_3099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3101 = 8'h1d == io_data_in[111:104] ? 8'ha4 : _GEN_3100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3102 = 8'h1e == io_data_in[111:104] ? 8'h72 : _GEN_3101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3103 = 8'h1f == io_data_in[111:104] ? 8'hc0 : _GEN_3102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3104 = 8'h20 == io_data_in[111:104] ? 8'hb7 : _GEN_3103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3105 = 8'h21 == io_data_in[111:104] ? 8'hfd : _GEN_3104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3106 = 8'h22 == io_data_in[111:104] ? 8'h93 : _GEN_3105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3107 = 8'h23 == io_data_in[111:104] ? 8'h26 : _GEN_3106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3108 = 8'h24 == io_data_in[111:104] ? 8'h36 : _GEN_3107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3109 = 8'h25 == io_data_in[111:104] ? 8'h3f : _GEN_3108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3110 = 8'h26 == io_data_in[111:104] ? 8'hf7 : _GEN_3109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3111 = 8'h27 == io_data_in[111:104] ? 8'hcc : _GEN_3110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3112 = 8'h28 == io_data_in[111:104] ? 8'h34 : _GEN_3111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3113 = 8'h29 == io_data_in[111:104] ? 8'ha5 : _GEN_3112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3114 = 8'h2a == io_data_in[111:104] ? 8'he5 : _GEN_3113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3115 = 8'h2b == io_data_in[111:104] ? 8'hf1 : _GEN_3114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3116 = 8'h2c == io_data_in[111:104] ? 8'h71 : _GEN_3115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3117 = 8'h2d == io_data_in[111:104] ? 8'hd8 : _GEN_3116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3118 = 8'h2e == io_data_in[111:104] ? 8'h31 : _GEN_3117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3119 = 8'h2f == io_data_in[111:104] ? 8'h15 : _GEN_3118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3120 = 8'h30 == io_data_in[111:104] ? 8'h4 : _GEN_3119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3121 = 8'h31 == io_data_in[111:104] ? 8'hc7 : _GEN_3120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3122 = 8'h32 == io_data_in[111:104] ? 8'h23 : _GEN_3121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3123 = 8'h33 == io_data_in[111:104] ? 8'hc3 : _GEN_3122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3124 = 8'h34 == io_data_in[111:104] ? 8'h18 : _GEN_3123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3125 = 8'h35 == io_data_in[111:104] ? 8'h96 : _GEN_3124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3126 = 8'h36 == io_data_in[111:104] ? 8'h5 : _GEN_3125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3127 = 8'h37 == io_data_in[111:104] ? 8'h9a : _GEN_3126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3128 = 8'h38 == io_data_in[111:104] ? 8'h7 : _GEN_3127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3129 = 8'h39 == io_data_in[111:104] ? 8'h12 : _GEN_3128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3130 = 8'h3a == io_data_in[111:104] ? 8'h80 : _GEN_3129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3131 = 8'h3b == io_data_in[111:104] ? 8'he2 : _GEN_3130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3132 = 8'h3c == io_data_in[111:104] ? 8'heb : _GEN_3131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3133 = 8'h3d == io_data_in[111:104] ? 8'h27 : _GEN_3132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3134 = 8'h3e == io_data_in[111:104] ? 8'hb2 : _GEN_3133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3135 = 8'h3f == io_data_in[111:104] ? 8'h75 : _GEN_3134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3136 = 8'h40 == io_data_in[111:104] ? 8'h9 : _GEN_3135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3137 = 8'h41 == io_data_in[111:104] ? 8'h83 : _GEN_3136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3138 = 8'h42 == io_data_in[111:104] ? 8'h2c : _GEN_3137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3139 = 8'h43 == io_data_in[111:104] ? 8'h1a : _GEN_3138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3140 = 8'h44 == io_data_in[111:104] ? 8'h1b : _GEN_3139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3141 = 8'h45 == io_data_in[111:104] ? 8'h6e : _GEN_3140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3142 = 8'h46 == io_data_in[111:104] ? 8'h5a : _GEN_3141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3143 = 8'h47 == io_data_in[111:104] ? 8'ha0 : _GEN_3142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3144 = 8'h48 == io_data_in[111:104] ? 8'h52 : _GEN_3143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3145 = 8'h49 == io_data_in[111:104] ? 8'h3b : _GEN_3144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3146 = 8'h4a == io_data_in[111:104] ? 8'hd6 : _GEN_3145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3147 = 8'h4b == io_data_in[111:104] ? 8'hb3 : _GEN_3146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3148 = 8'h4c == io_data_in[111:104] ? 8'h29 : _GEN_3147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3149 = 8'h4d == io_data_in[111:104] ? 8'he3 : _GEN_3148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3150 = 8'h4e == io_data_in[111:104] ? 8'h2f : _GEN_3149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3151 = 8'h4f == io_data_in[111:104] ? 8'h84 : _GEN_3150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3152 = 8'h50 == io_data_in[111:104] ? 8'h53 : _GEN_3151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3153 = 8'h51 == io_data_in[111:104] ? 8'hd1 : _GEN_3152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3154 = 8'h52 == io_data_in[111:104] ? 8'h0 : _GEN_3153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3155 = 8'h53 == io_data_in[111:104] ? 8'hed : _GEN_3154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3156 = 8'h54 == io_data_in[111:104] ? 8'h20 : _GEN_3155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3157 = 8'h55 == io_data_in[111:104] ? 8'hfc : _GEN_3156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3158 = 8'h56 == io_data_in[111:104] ? 8'hb1 : _GEN_3157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3159 = 8'h57 == io_data_in[111:104] ? 8'h5b : _GEN_3158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3160 = 8'h58 == io_data_in[111:104] ? 8'h6a : _GEN_3159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3161 = 8'h59 == io_data_in[111:104] ? 8'hcb : _GEN_3160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3162 = 8'h5a == io_data_in[111:104] ? 8'hbe : _GEN_3161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3163 = 8'h5b == io_data_in[111:104] ? 8'h39 : _GEN_3162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3164 = 8'h5c == io_data_in[111:104] ? 8'h4a : _GEN_3163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3165 = 8'h5d == io_data_in[111:104] ? 8'h4c : _GEN_3164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3166 = 8'h5e == io_data_in[111:104] ? 8'h58 : _GEN_3165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3167 = 8'h5f == io_data_in[111:104] ? 8'hcf : _GEN_3166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3168 = 8'h60 == io_data_in[111:104] ? 8'hd0 : _GEN_3167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3169 = 8'h61 == io_data_in[111:104] ? 8'hef : _GEN_3168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3170 = 8'h62 == io_data_in[111:104] ? 8'haa : _GEN_3169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3171 = 8'h63 == io_data_in[111:104] ? 8'hfb : _GEN_3170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3172 = 8'h64 == io_data_in[111:104] ? 8'h43 : _GEN_3171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3173 = 8'h65 == io_data_in[111:104] ? 8'h4d : _GEN_3172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3174 = 8'h66 == io_data_in[111:104] ? 8'h33 : _GEN_3173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3175 = 8'h67 == io_data_in[111:104] ? 8'h85 : _GEN_3174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3176 = 8'h68 == io_data_in[111:104] ? 8'h45 : _GEN_3175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3177 = 8'h69 == io_data_in[111:104] ? 8'hf9 : _GEN_3176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3178 = 8'h6a == io_data_in[111:104] ? 8'h2 : _GEN_3177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3179 = 8'h6b == io_data_in[111:104] ? 8'h7f : _GEN_3178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3180 = 8'h6c == io_data_in[111:104] ? 8'h50 : _GEN_3179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3181 = 8'h6d == io_data_in[111:104] ? 8'h3c : _GEN_3180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3182 = 8'h6e == io_data_in[111:104] ? 8'h9f : _GEN_3181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3183 = 8'h6f == io_data_in[111:104] ? 8'ha8 : _GEN_3182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3184 = 8'h70 == io_data_in[111:104] ? 8'h51 : _GEN_3183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3185 = 8'h71 == io_data_in[111:104] ? 8'ha3 : _GEN_3184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3186 = 8'h72 == io_data_in[111:104] ? 8'h40 : _GEN_3185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3187 = 8'h73 == io_data_in[111:104] ? 8'h8f : _GEN_3186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3188 = 8'h74 == io_data_in[111:104] ? 8'h92 : _GEN_3187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3189 = 8'h75 == io_data_in[111:104] ? 8'h9d : _GEN_3188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3190 = 8'h76 == io_data_in[111:104] ? 8'h38 : _GEN_3189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3191 = 8'h77 == io_data_in[111:104] ? 8'hf5 : _GEN_3190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3192 = 8'h78 == io_data_in[111:104] ? 8'hbc : _GEN_3191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3193 = 8'h79 == io_data_in[111:104] ? 8'hb6 : _GEN_3192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3194 = 8'h7a == io_data_in[111:104] ? 8'hda : _GEN_3193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3195 = 8'h7b == io_data_in[111:104] ? 8'h21 : _GEN_3194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3196 = 8'h7c == io_data_in[111:104] ? 8'h10 : _GEN_3195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3197 = 8'h7d == io_data_in[111:104] ? 8'hff : _GEN_3196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3198 = 8'h7e == io_data_in[111:104] ? 8'hf3 : _GEN_3197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3199 = 8'h7f == io_data_in[111:104] ? 8'hd2 : _GEN_3198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3200 = 8'h80 == io_data_in[111:104] ? 8'hcd : _GEN_3199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3201 = 8'h81 == io_data_in[111:104] ? 8'hc : _GEN_3200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3202 = 8'h82 == io_data_in[111:104] ? 8'h13 : _GEN_3201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3203 = 8'h83 == io_data_in[111:104] ? 8'hec : _GEN_3202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3204 = 8'h84 == io_data_in[111:104] ? 8'h5f : _GEN_3203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3205 = 8'h85 == io_data_in[111:104] ? 8'h97 : _GEN_3204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3206 = 8'h86 == io_data_in[111:104] ? 8'h44 : _GEN_3205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3207 = 8'h87 == io_data_in[111:104] ? 8'h17 : _GEN_3206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3208 = 8'h88 == io_data_in[111:104] ? 8'hc4 : _GEN_3207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3209 = 8'h89 == io_data_in[111:104] ? 8'ha7 : _GEN_3208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3210 = 8'h8a == io_data_in[111:104] ? 8'h7e : _GEN_3209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3211 = 8'h8b == io_data_in[111:104] ? 8'h3d : _GEN_3210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3212 = 8'h8c == io_data_in[111:104] ? 8'h64 : _GEN_3211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3213 = 8'h8d == io_data_in[111:104] ? 8'h5d : _GEN_3212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3214 = 8'h8e == io_data_in[111:104] ? 8'h19 : _GEN_3213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3215 = 8'h8f == io_data_in[111:104] ? 8'h73 : _GEN_3214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3216 = 8'h90 == io_data_in[111:104] ? 8'h60 : _GEN_3215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3217 = 8'h91 == io_data_in[111:104] ? 8'h81 : _GEN_3216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3218 = 8'h92 == io_data_in[111:104] ? 8'h4f : _GEN_3217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3219 = 8'h93 == io_data_in[111:104] ? 8'hdc : _GEN_3218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3220 = 8'h94 == io_data_in[111:104] ? 8'h22 : _GEN_3219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3221 = 8'h95 == io_data_in[111:104] ? 8'h2a : _GEN_3220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3222 = 8'h96 == io_data_in[111:104] ? 8'h90 : _GEN_3221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3223 = 8'h97 == io_data_in[111:104] ? 8'h88 : _GEN_3222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3224 = 8'h98 == io_data_in[111:104] ? 8'h46 : _GEN_3223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3225 = 8'h99 == io_data_in[111:104] ? 8'hee : _GEN_3224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3226 = 8'h9a == io_data_in[111:104] ? 8'hb8 : _GEN_3225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3227 = 8'h9b == io_data_in[111:104] ? 8'h14 : _GEN_3226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3228 = 8'h9c == io_data_in[111:104] ? 8'hde : _GEN_3227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3229 = 8'h9d == io_data_in[111:104] ? 8'h5e : _GEN_3228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3230 = 8'h9e == io_data_in[111:104] ? 8'hb : _GEN_3229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3231 = 8'h9f == io_data_in[111:104] ? 8'hdb : _GEN_3230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3232 = 8'ha0 == io_data_in[111:104] ? 8'he0 : _GEN_3231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3233 = 8'ha1 == io_data_in[111:104] ? 8'h32 : _GEN_3232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3234 = 8'ha2 == io_data_in[111:104] ? 8'h3a : _GEN_3233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3235 = 8'ha3 == io_data_in[111:104] ? 8'ha : _GEN_3234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3236 = 8'ha4 == io_data_in[111:104] ? 8'h49 : _GEN_3235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3237 = 8'ha5 == io_data_in[111:104] ? 8'h6 : _GEN_3236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3238 = 8'ha6 == io_data_in[111:104] ? 8'h24 : _GEN_3237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3239 = 8'ha7 == io_data_in[111:104] ? 8'h5c : _GEN_3238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3240 = 8'ha8 == io_data_in[111:104] ? 8'hc2 : _GEN_3239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3241 = 8'ha9 == io_data_in[111:104] ? 8'hd3 : _GEN_3240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3242 = 8'haa == io_data_in[111:104] ? 8'hac : _GEN_3241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3243 = 8'hab == io_data_in[111:104] ? 8'h62 : _GEN_3242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3244 = 8'hac == io_data_in[111:104] ? 8'h91 : _GEN_3243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3245 = 8'had == io_data_in[111:104] ? 8'h95 : _GEN_3244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3246 = 8'hae == io_data_in[111:104] ? 8'he4 : _GEN_3245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3247 = 8'haf == io_data_in[111:104] ? 8'h79 : _GEN_3246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3248 = 8'hb0 == io_data_in[111:104] ? 8'he7 : _GEN_3247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3249 = 8'hb1 == io_data_in[111:104] ? 8'hc8 : _GEN_3248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3250 = 8'hb2 == io_data_in[111:104] ? 8'h37 : _GEN_3249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3251 = 8'hb3 == io_data_in[111:104] ? 8'h6d : _GEN_3250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3252 = 8'hb4 == io_data_in[111:104] ? 8'h8d : _GEN_3251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3253 = 8'hb5 == io_data_in[111:104] ? 8'hd5 : _GEN_3252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3254 = 8'hb6 == io_data_in[111:104] ? 8'h4e : _GEN_3253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3255 = 8'hb7 == io_data_in[111:104] ? 8'ha9 : _GEN_3254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3256 = 8'hb8 == io_data_in[111:104] ? 8'h6c : _GEN_3255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3257 = 8'hb9 == io_data_in[111:104] ? 8'h56 : _GEN_3256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3258 = 8'hba == io_data_in[111:104] ? 8'hf4 : _GEN_3257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3259 = 8'hbb == io_data_in[111:104] ? 8'hea : _GEN_3258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3260 = 8'hbc == io_data_in[111:104] ? 8'h65 : _GEN_3259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3261 = 8'hbd == io_data_in[111:104] ? 8'h7a : _GEN_3260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3262 = 8'hbe == io_data_in[111:104] ? 8'hae : _GEN_3261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3263 = 8'hbf == io_data_in[111:104] ? 8'h8 : _GEN_3262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3264 = 8'hc0 == io_data_in[111:104] ? 8'hba : _GEN_3263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3265 = 8'hc1 == io_data_in[111:104] ? 8'h78 : _GEN_3264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3266 = 8'hc2 == io_data_in[111:104] ? 8'h25 : _GEN_3265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3267 = 8'hc3 == io_data_in[111:104] ? 8'h2e : _GEN_3266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3268 = 8'hc4 == io_data_in[111:104] ? 8'h1c : _GEN_3267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3269 = 8'hc5 == io_data_in[111:104] ? 8'ha6 : _GEN_3268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3270 = 8'hc6 == io_data_in[111:104] ? 8'hb4 : _GEN_3269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3271 = 8'hc7 == io_data_in[111:104] ? 8'hc6 : _GEN_3270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3272 = 8'hc8 == io_data_in[111:104] ? 8'he8 : _GEN_3271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3273 = 8'hc9 == io_data_in[111:104] ? 8'hdd : _GEN_3272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3274 = 8'hca == io_data_in[111:104] ? 8'h74 : _GEN_3273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3275 = 8'hcb == io_data_in[111:104] ? 8'h1f : _GEN_3274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3276 = 8'hcc == io_data_in[111:104] ? 8'h4b : _GEN_3275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3277 = 8'hcd == io_data_in[111:104] ? 8'hbd : _GEN_3276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3278 = 8'hce == io_data_in[111:104] ? 8'h8b : _GEN_3277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3279 = 8'hcf == io_data_in[111:104] ? 8'h8a : _GEN_3278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3280 = 8'hd0 == io_data_in[111:104] ? 8'h70 : _GEN_3279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3281 = 8'hd1 == io_data_in[111:104] ? 8'h3e : _GEN_3280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3282 = 8'hd2 == io_data_in[111:104] ? 8'hb5 : _GEN_3281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3283 = 8'hd3 == io_data_in[111:104] ? 8'h66 : _GEN_3282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3284 = 8'hd4 == io_data_in[111:104] ? 8'h48 : _GEN_3283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3285 = 8'hd5 == io_data_in[111:104] ? 8'h3 : _GEN_3284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3286 = 8'hd6 == io_data_in[111:104] ? 8'hf6 : _GEN_3285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3287 = 8'hd7 == io_data_in[111:104] ? 8'he : _GEN_3286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3288 = 8'hd8 == io_data_in[111:104] ? 8'h61 : _GEN_3287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3289 = 8'hd9 == io_data_in[111:104] ? 8'h35 : _GEN_3288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3290 = 8'hda == io_data_in[111:104] ? 8'h57 : _GEN_3289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3291 = 8'hdb == io_data_in[111:104] ? 8'hb9 : _GEN_3290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3292 = 8'hdc == io_data_in[111:104] ? 8'h86 : _GEN_3291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3293 = 8'hdd == io_data_in[111:104] ? 8'hc1 : _GEN_3292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3294 = 8'hde == io_data_in[111:104] ? 8'h1d : _GEN_3293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3295 = 8'hdf == io_data_in[111:104] ? 8'h9e : _GEN_3294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3296 = 8'he0 == io_data_in[111:104] ? 8'he1 : _GEN_3295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3297 = 8'he1 == io_data_in[111:104] ? 8'hf8 : _GEN_3296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3298 = 8'he2 == io_data_in[111:104] ? 8'h98 : _GEN_3297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3299 = 8'he3 == io_data_in[111:104] ? 8'h11 : _GEN_3298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3300 = 8'he4 == io_data_in[111:104] ? 8'h69 : _GEN_3299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3301 = 8'he5 == io_data_in[111:104] ? 8'hd9 : _GEN_3300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3302 = 8'he6 == io_data_in[111:104] ? 8'h8e : _GEN_3301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3303 = 8'he7 == io_data_in[111:104] ? 8'h94 : _GEN_3302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3304 = 8'he8 == io_data_in[111:104] ? 8'h9b : _GEN_3303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3305 = 8'he9 == io_data_in[111:104] ? 8'h1e : _GEN_3304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3306 = 8'hea == io_data_in[111:104] ? 8'h87 : _GEN_3305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3307 = 8'heb == io_data_in[111:104] ? 8'he9 : _GEN_3306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3308 = 8'hec == io_data_in[111:104] ? 8'hce : _GEN_3307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3309 = 8'hed == io_data_in[111:104] ? 8'h55 : _GEN_3308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3310 = 8'hee == io_data_in[111:104] ? 8'h28 : _GEN_3309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3311 = 8'hef == io_data_in[111:104] ? 8'hdf : _GEN_3310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3312 = 8'hf0 == io_data_in[111:104] ? 8'h8c : _GEN_3311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3313 = 8'hf1 == io_data_in[111:104] ? 8'ha1 : _GEN_3312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3314 = 8'hf2 == io_data_in[111:104] ? 8'h89 : _GEN_3313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3315 = 8'hf3 == io_data_in[111:104] ? 8'hd : _GEN_3314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3316 = 8'hf4 == io_data_in[111:104] ? 8'hbf : _GEN_3315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3317 = 8'hf5 == io_data_in[111:104] ? 8'he6 : _GEN_3316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3318 = 8'hf6 == io_data_in[111:104] ? 8'h42 : _GEN_3317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3319 = 8'hf7 == io_data_in[111:104] ? 8'h68 : _GEN_3318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3320 = 8'hf8 == io_data_in[111:104] ? 8'h41 : _GEN_3319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3321 = 8'hf9 == io_data_in[111:104] ? 8'h99 : _GEN_3320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3322 = 8'hfa == io_data_in[111:104] ? 8'h2d : _GEN_3321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3323 = 8'hfb == io_data_in[111:104] ? 8'hf : _GEN_3322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3324 = 8'hfc == io_data_in[111:104] ? 8'hb0 : _GEN_3323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3325 = 8'hfd == io_data_in[111:104] ? 8'h54 : _GEN_3324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3326 = 8'hfe == io_data_in[111:104] ? 8'hbb : _GEN_3325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3327 = 8'hff == io_data_in[111:104] ? 8'h16 : _GEN_3326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3329 = 8'h1 == io_data_in[103:96] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3330 = 8'h2 == io_data_in[103:96] ? 8'h77 : _GEN_3329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3331 = 8'h3 == io_data_in[103:96] ? 8'h7b : _GEN_3330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3332 = 8'h4 == io_data_in[103:96] ? 8'hf2 : _GEN_3331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3333 = 8'h5 == io_data_in[103:96] ? 8'h6b : _GEN_3332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3334 = 8'h6 == io_data_in[103:96] ? 8'h6f : _GEN_3333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3335 = 8'h7 == io_data_in[103:96] ? 8'hc5 : _GEN_3334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3336 = 8'h8 == io_data_in[103:96] ? 8'h30 : _GEN_3335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3337 = 8'h9 == io_data_in[103:96] ? 8'h1 : _GEN_3336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3338 = 8'ha == io_data_in[103:96] ? 8'h67 : _GEN_3337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3339 = 8'hb == io_data_in[103:96] ? 8'h2b : _GEN_3338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3340 = 8'hc == io_data_in[103:96] ? 8'hfe : _GEN_3339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3341 = 8'hd == io_data_in[103:96] ? 8'hd7 : _GEN_3340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3342 = 8'he == io_data_in[103:96] ? 8'hab : _GEN_3341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3343 = 8'hf == io_data_in[103:96] ? 8'h76 : _GEN_3342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3344 = 8'h10 == io_data_in[103:96] ? 8'hca : _GEN_3343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3345 = 8'h11 == io_data_in[103:96] ? 8'h82 : _GEN_3344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3346 = 8'h12 == io_data_in[103:96] ? 8'hc9 : _GEN_3345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3347 = 8'h13 == io_data_in[103:96] ? 8'h7d : _GEN_3346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3348 = 8'h14 == io_data_in[103:96] ? 8'hfa : _GEN_3347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3349 = 8'h15 == io_data_in[103:96] ? 8'h59 : _GEN_3348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3350 = 8'h16 == io_data_in[103:96] ? 8'h47 : _GEN_3349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3351 = 8'h17 == io_data_in[103:96] ? 8'hf0 : _GEN_3350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3352 = 8'h18 == io_data_in[103:96] ? 8'had : _GEN_3351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3353 = 8'h19 == io_data_in[103:96] ? 8'hd4 : _GEN_3352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3354 = 8'h1a == io_data_in[103:96] ? 8'ha2 : _GEN_3353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3355 = 8'h1b == io_data_in[103:96] ? 8'haf : _GEN_3354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3356 = 8'h1c == io_data_in[103:96] ? 8'h9c : _GEN_3355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3357 = 8'h1d == io_data_in[103:96] ? 8'ha4 : _GEN_3356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3358 = 8'h1e == io_data_in[103:96] ? 8'h72 : _GEN_3357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3359 = 8'h1f == io_data_in[103:96] ? 8'hc0 : _GEN_3358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3360 = 8'h20 == io_data_in[103:96] ? 8'hb7 : _GEN_3359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3361 = 8'h21 == io_data_in[103:96] ? 8'hfd : _GEN_3360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3362 = 8'h22 == io_data_in[103:96] ? 8'h93 : _GEN_3361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3363 = 8'h23 == io_data_in[103:96] ? 8'h26 : _GEN_3362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3364 = 8'h24 == io_data_in[103:96] ? 8'h36 : _GEN_3363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3365 = 8'h25 == io_data_in[103:96] ? 8'h3f : _GEN_3364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3366 = 8'h26 == io_data_in[103:96] ? 8'hf7 : _GEN_3365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3367 = 8'h27 == io_data_in[103:96] ? 8'hcc : _GEN_3366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3368 = 8'h28 == io_data_in[103:96] ? 8'h34 : _GEN_3367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3369 = 8'h29 == io_data_in[103:96] ? 8'ha5 : _GEN_3368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3370 = 8'h2a == io_data_in[103:96] ? 8'he5 : _GEN_3369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3371 = 8'h2b == io_data_in[103:96] ? 8'hf1 : _GEN_3370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3372 = 8'h2c == io_data_in[103:96] ? 8'h71 : _GEN_3371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3373 = 8'h2d == io_data_in[103:96] ? 8'hd8 : _GEN_3372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3374 = 8'h2e == io_data_in[103:96] ? 8'h31 : _GEN_3373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3375 = 8'h2f == io_data_in[103:96] ? 8'h15 : _GEN_3374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3376 = 8'h30 == io_data_in[103:96] ? 8'h4 : _GEN_3375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3377 = 8'h31 == io_data_in[103:96] ? 8'hc7 : _GEN_3376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3378 = 8'h32 == io_data_in[103:96] ? 8'h23 : _GEN_3377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3379 = 8'h33 == io_data_in[103:96] ? 8'hc3 : _GEN_3378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3380 = 8'h34 == io_data_in[103:96] ? 8'h18 : _GEN_3379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3381 = 8'h35 == io_data_in[103:96] ? 8'h96 : _GEN_3380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3382 = 8'h36 == io_data_in[103:96] ? 8'h5 : _GEN_3381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3383 = 8'h37 == io_data_in[103:96] ? 8'h9a : _GEN_3382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3384 = 8'h38 == io_data_in[103:96] ? 8'h7 : _GEN_3383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3385 = 8'h39 == io_data_in[103:96] ? 8'h12 : _GEN_3384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3386 = 8'h3a == io_data_in[103:96] ? 8'h80 : _GEN_3385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3387 = 8'h3b == io_data_in[103:96] ? 8'he2 : _GEN_3386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3388 = 8'h3c == io_data_in[103:96] ? 8'heb : _GEN_3387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3389 = 8'h3d == io_data_in[103:96] ? 8'h27 : _GEN_3388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3390 = 8'h3e == io_data_in[103:96] ? 8'hb2 : _GEN_3389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3391 = 8'h3f == io_data_in[103:96] ? 8'h75 : _GEN_3390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3392 = 8'h40 == io_data_in[103:96] ? 8'h9 : _GEN_3391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3393 = 8'h41 == io_data_in[103:96] ? 8'h83 : _GEN_3392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3394 = 8'h42 == io_data_in[103:96] ? 8'h2c : _GEN_3393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3395 = 8'h43 == io_data_in[103:96] ? 8'h1a : _GEN_3394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3396 = 8'h44 == io_data_in[103:96] ? 8'h1b : _GEN_3395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3397 = 8'h45 == io_data_in[103:96] ? 8'h6e : _GEN_3396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3398 = 8'h46 == io_data_in[103:96] ? 8'h5a : _GEN_3397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3399 = 8'h47 == io_data_in[103:96] ? 8'ha0 : _GEN_3398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3400 = 8'h48 == io_data_in[103:96] ? 8'h52 : _GEN_3399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3401 = 8'h49 == io_data_in[103:96] ? 8'h3b : _GEN_3400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3402 = 8'h4a == io_data_in[103:96] ? 8'hd6 : _GEN_3401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3403 = 8'h4b == io_data_in[103:96] ? 8'hb3 : _GEN_3402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3404 = 8'h4c == io_data_in[103:96] ? 8'h29 : _GEN_3403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3405 = 8'h4d == io_data_in[103:96] ? 8'he3 : _GEN_3404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3406 = 8'h4e == io_data_in[103:96] ? 8'h2f : _GEN_3405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3407 = 8'h4f == io_data_in[103:96] ? 8'h84 : _GEN_3406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3408 = 8'h50 == io_data_in[103:96] ? 8'h53 : _GEN_3407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3409 = 8'h51 == io_data_in[103:96] ? 8'hd1 : _GEN_3408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3410 = 8'h52 == io_data_in[103:96] ? 8'h0 : _GEN_3409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3411 = 8'h53 == io_data_in[103:96] ? 8'hed : _GEN_3410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3412 = 8'h54 == io_data_in[103:96] ? 8'h20 : _GEN_3411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3413 = 8'h55 == io_data_in[103:96] ? 8'hfc : _GEN_3412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3414 = 8'h56 == io_data_in[103:96] ? 8'hb1 : _GEN_3413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3415 = 8'h57 == io_data_in[103:96] ? 8'h5b : _GEN_3414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3416 = 8'h58 == io_data_in[103:96] ? 8'h6a : _GEN_3415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3417 = 8'h59 == io_data_in[103:96] ? 8'hcb : _GEN_3416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3418 = 8'h5a == io_data_in[103:96] ? 8'hbe : _GEN_3417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3419 = 8'h5b == io_data_in[103:96] ? 8'h39 : _GEN_3418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3420 = 8'h5c == io_data_in[103:96] ? 8'h4a : _GEN_3419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3421 = 8'h5d == io_data_in[103:96] ? 8'h4c : _GEN_3420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3422 = 8'h5e == io_data_in[103:96] ? 8'h58 : _GEN_3421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3423 = 8'h5f == io_data_in[103:96] ? 8'hcf : _GEN_3422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3424 = 8'h60 == io_data_in[103:96] ? 8'hd0 : _GEN_3423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3425 = 8'h61 == io_data_in[103:96] ? 8'hef : _GEN_3424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3426 = 8'h62 == io_data_in[103:96] ? 8'haa : _GEN_3425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3427 = 8'h63 == io_data_in[103:96] ? 8'hfb : _GEN_3426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3428 = 8'h64 == io_data_in[103:96] ? 8'h43 : _GEN_3427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3429 = 8'h65 == io_data_in[103:96] ? 8'h4d : _GEN_3428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3430 = 8'h66 == io_data_in[103:96] ? 8'h33 : _GEN_3429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3431 = 8'h67 == io_data_in[103:96] ? 8'h85 : _GEN_3430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3432 = 8'h68 == io_data_in[103:96] ? 8'h45 : _GEN_3431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3433 = 8'h69 == io_data_in[103:96] ? 8'hf9 : _GEN_3432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3434 = 8'h6a == io_data_in[103:96] ? 8'h2 : _GEN_3433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3435 = 8'h6b == io_data_in[103:96] ? 8'h7f : _GEN_3434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3436 = 8'h6c == io_data_in[103:96] ? 8'h50 : _GEN_3435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3437 = 8'h6d == io_data_in[103:96] ? 8'h3c : _GEN_3436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3438 = 8'h6e == io_data_in[103:96] ? 8'h9f : _GEN_3437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3439 = 8'h6f == io_data_in[103:96] ? 8'ha8 : _GEN_3438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3440 = 8'h70 == io_data_in[103:96] ? 8'h51 : _GEN_3439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3441 = 8'h71 == io_data_in[103:96] ? 8'ha3 : _GEN_3440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3442 = 8'h72 == io_data_in[103:96] ? 8'h40 : _GEN_3441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3443 = 8'h73 == io_data_in[103:96] ? 8'h8f : _GEN_3442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3444 = 8'h74 == io_data_in[103:96] ? 8'h92 : _GEN_3443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3445 = 8'h75 == io_data_in[103:96] ? 8'h9d : _GEN_3444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3446 = 8'h76 == io_data_in[103:96] ? 8'h38 : _GEN_3445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3447 = 8'h77 == io_data_in[103:96] ? 8'hf5 : _GEN_3446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3448 = 8'h78 == io_data_in[103:96] ? 8'hbc : _GEN_3447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3449 = 8'h79 == io_data_in[103:96] ? 8'hb6 : _GEN_3448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3450 = 8'h7a == io_data_in[103:96] ? 8'hda : _GEN_3449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3451 = 8'h7b == io_data_in[103:96] ? 8'h21 : _GEN_3450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3452 = 8'h7c == io_data_in[103:96] ? 8'h10 : _GEN_3451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3453 = 8'h7d == io_data_in[103:96] ? 8'hff : _GEN_3452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3454 = 8'h7e == io_data_in[103:96] ? 8'hf3 : _GEN_3453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3455 = 8'h7f == io_data_in[103:96] ? 8'hd2 : _GEN_3454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3456 = 8'h80 == io_data_in[103:96] ? 8'hcd : _GEN_3455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3457 = 8'h81 == io_data_in[103:96] ? 8'hc : _GEN_3456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3458 = 8'h82 == io_data_in[103:96] ? 8'h13 : _GEN_3457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3459 = 8'h83 == io_data_in[103:96] ? 8'hec : _GEN_3458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3460 = 8'h84 == io_data_in[103:96] ? 8'h5f : _GEN_3459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3461 = 8'h85 == io_data_in[103:96] ? 8'h97 : _GEN_3460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3462 = 8'h86 == io_data_in[103:96] ? 8'h44 : _GEN_3461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3463 = 8'h87 == io_data_in[103:96] ? 8'h17 : _GEN_3462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3464 = 8'h88 == io_data_in[103:96] ? 8'hc4 : _GEN_3463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3465 = 8'h89 == io_data_in[103:96] ? 8'ha7 : _GEN_3464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3466 = 8'h8a == io_data_in[103:96] ? 8'h7e : _GEN_3465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3467 = 8'h8b == io_data_in[103:96] ? 8'h3d : _GEN_3466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3468 = 8'h8c == io_data_in[103:96] ? 8'h64 : _GEN_3467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3469 = 8'h8d == io_data_in[103:96] ? 8'h5d : _GEN_3468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3470 = 8'h8e == io_data_in[103:96] ? 8'h19 : _GEN_3469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3471 = 8'h8f == io_data_in[103:96] ? 8'h73 : _GEN_3470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3472 = 8'h90 == io_data_in[103:96] ? 8'h60 : _GEN_3471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3473 = 8'h91 == io_data_in[103:96] ? 8'h81 : _GEN_3472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3474 = 8'h92 == io_data_in[103:96] ? 8'h4f : _GEN_3473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3475 = 8'h93 == io_data_in[103:96] ? 8'hdc : _GEN_3474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3476 = 8'h94 == io_data_in[103:96] ? 8'h22 : _GEN_3475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3477 = 8'h95 == io_data_in[103:96] ? 8'h2a : _GEN_3476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3478 = 8'h96 == io_data_in[103:96] ? 8'h90 : _GEN_3477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3479 = 8'h97 == io_data_in[103:96] ? 8'h88 : _GEN_3478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3480 = 8'h98 == io_data_in[103:96] ? 8'h46 : _GEN_3479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3481 = 8'h99 == io_data_in[103:96] ? 8'hee : _GEN_3480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3482 = 8'h9a == io_data_in[103:96] ? 8'hb8 : _GEN_3481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3483 = 8'h9b == io_data_in[103:96] ? 8'h14 : _GEN_3482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3484 = 8'h9c == io_data_in[103:96] ? 8'hde : _GEN_3483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3485 = 8'h9d == io_data_in[103:96] ? 8'h5e : _GEN_3484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3486 = 8'h9e == io_data_in[103:96] ? 8'hb : _GEN_3485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3487 = 8'h9f == io_data_in[103:96] ? 8'hdb : _GEN_3486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3488 = 8'ha0 == io_data_in[103:96] ? 8'he0 : _GEN_3487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3489 = 8'ha1 == io_data_in[103:96] ? 8'h32 : _GEN_3488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3490 = 8'ha2 == io_data_in[103:96] ? 8'h3a : _GEN_3489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3491 = 8'ha3 == io_data_in[103:96] ? 8'ha : _GEN_3490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3492 = 8'ha4 == io_data_in[103:96] ? 8'h49 : _GEN_3491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3493 = 8'ha5 == io_data_in[103:96] ? 8'h6 : _GEN_3492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3494 = 8'ha6 == io_data_in[103:96] ? 8'h24 : _GEN_3493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3495 = 8'ha7 == io_data_in[103:96] ? 8'h5c : _GEN_3494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3496 = 8'ha8 == io_data_in[103:96] ? 8'hc2 : _GEN_3495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3497 = 8'ha9 == io_data_in[103:96] ? 8'hd3 : _GEN_3496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3498 = 8'haa == io_data_in[103:96] ? 8'hac : _GEN_3497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3499 = 8'hab == io_data_in[103:96] ? 8'h62 : _GEN_3498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3500 = 8'hac == io_data_in[103:96] ? 8'h91 : _GEN_3499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3501 = 8'had == io_data_in[103:96] ? 8'h95 : _GEN_3500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3502 = 8'hae == io_data_in[103:96] ? 8'he4 : _GEN_3501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3503 = 8'haf == io_data_in[103:96] ? 8'h79 : _GEN_3502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3504 = 8'hb0 == io_data_in[103:96] ? 8'he7 : _GEN_3503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3505 = 8'hb1 == io_data_in[103:96] ? 8'hc8 : _GEN_3504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3506 = 8'hb2 == io_data_in[103:96] ? 8'h37 : _GEN_3505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3507 = 8'hb3 == io_data_in[103:96] ? 8'h6d : _GEN_3506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3508 = 8'hb4 == io_data_in[103:96] ? 8'h8d : _GEN_3507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3509 = 8'hb5 == io_data_in[103:96] ? 8'hd5 : _GEN_3508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3510 = 8'hb6 == io_data_in[103:96] ? 8'h4e : _GEN_3509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3511 = 8'hb7 == io_data_in[103:96] ? 8'ha9 : _GEN_3510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3512 = 8'hb8 == io_data_in[103:96] ? 8'h6c : _GEN_3511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3513 = 8'hb9 == io_data_in[103:96] ? 8'h56 : _GEN_3512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3514 = 8'hba == io_data_in[103:96] ? 8'hf4 : _GEN_3513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3515 = 8'hbb == io_data_in[103:96] ? 8'hea : _GEN_3514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3516 = 8'hbc == io_data_in[103:96] ? 8'h65 : _GEN_3515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3517 = 8'hbd == io_data_in[103:96] ? 8'h7a : _GEN_3516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3518 = 8'hbe == io_data_in[103:96] ? 8'hae : _GEN_3517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3519 = 8'hbf == io_data_in[103:96] ? 8'h8 : _GEN_3518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3520 = 8'hc0 == io_data_in[103:96] ? 8'hba : _GEN_3519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3521 = 8'hc1 == io_data_in[103:96] ? 8'h78 : _GEN_3520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3522 = 8'hc2 == io_data_in[103:96] ? 8'h25 : _GEN_3521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3523 = 8'hc3 == io_data_in[103:96] ? 8'h2e : _GEN_3522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3524 = 8'hc4 == io_data_in[103:96] ? 8'h1c : _GEN_3523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3525 = 8'hc5 == io_data_in[103:96] ? 8'ha6 : _GEN_3524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3526 = 8'hc6 == io_data_in[103:96] ? 8'hb4 : _GEN_3525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3527 = 8'hc7 == io_data_in[103:96] ? 8'hc6 : _GEN_3526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3528 = 8'hc8 == io_data_in[103:96] ? 8'he8 : _GEN_3527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3529 = 8'hc9 == io_data_in[103:96] ? 8'hdd : _GEN_3528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3530 = 8'hca == io_data_in[103:96] ? 8'h74 : _GEN_3529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3531 = 8'hcb == io_data_in[103:96] ? 8'h1f : _GEN_3530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3532 = 8'hcc == io_data_in[103:96] ? 8'h4b : _GEN_3531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3533 = 8'hcd == io_data_in[103:96] ? 8'hbd : _GEN_3532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3534 = 8'hce == io_data_in[103:96] ? 8'h8b : _GEN_3533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3535 = 8'hcf == io_data_in[103:96] ? 8'h8a : _GEN_3534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3536 = 8'hd0 == io_data_in[103:96] ? 8'h70 : _GEN_3535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3537 = 8'hd1 == io_data_in[103:96] ? 8'h3e : _GEN_3536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3538 = 8'hd2 == io_data_in[103:96] ? 8'hb5 : _GEN_3537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3539 = 8'hd3 == io_data_in[103:96] ? 8'h66 : _GEN_3538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3540 = 8'hd4 == io_data_in[103:96] ? 8'h48 : _GEN_3539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3541 = 8'hd5 == io_data_in[103:96] ? 8'h3 : _GEN_3540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3542 = 8'hd6 == io_data_in[103:96] ? 8'hf6 : _GEN_3541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3543 = 8'hd7 == io_data_in[103:96] ? 8'he : _GEN_3542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3544 = 8'hd8 == io_data_in[103:96] ? 8'h61 : _GEN_3543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3545 = 8'hd9 == io_data_in[103:96] ? 8'h35 : _GEN_3544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3546 = 8'hda == io_data_in[103:96] ? 8'h57 : _GEN_3545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3547 = 8'hdb == io_data_in[103:96] ? 8'hb9 : _GEN_3546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3548 = 8'hdc == io_data_in[103:96] ? 8'h86 : _GEN_3547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3549 = 8'hdd == io_data_in[103:96] ? 8'hc1 : _GEN_3548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3550 = 8'hde == io_data_in[103:96] ? 8'h1d : _GEN_3549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3551 = 8'hdf == io_data_in[103:96] ? 8'h9e : _GEN_3550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3552 = 8'he0 == io_data_in[103:96] ? 8'he1 : _GEN_3551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3553 = 8'he1 == io_data_in[103:96] ? 8'hf8 : _GEN_3552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3554 = 8'he2 == io_data_in[103:96] ? 8'h98 : _GEN_3553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3555 = 8'he3 == io_data_in[103:96] ? 8'h11 : _GEN_3554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3556 = 8'he4 == io_data_in[103:96] ? 8'h69 : _GEN_3555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3557 = 8'he5 == io_data_in[103:96] ? 8'hd9 : _GEN_3556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3558 = 8'he6 == io_data_in[103:96] ? 8'h8e : _GEN_3557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3559 = 8'he7 == io_data_in[103:96] ? 8'h94 : _GEN_3558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3560 = 8'he8 == io_data_in[103:96] ? 8'h9b : _GEN_3559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3561 = 8'he9 == io_data_in[103:96] ? 8'h1e : _GEN_3560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3562 = 8'hea == io_data_in[103:96] ? 8'h87 : _GEN_3561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3563 = 8'heb == io_data_in[103:96] ? 8'he9 : _GEN_3562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3564 = 8'hec == io_data_in[103:96] ? 8'hce : _GEN_3563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3565 = 8'hed == io_data_in[103:96] ? 8'h55 : _GEN_3564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3566 = 8'hee == io_data_in[103:96] ? 8'h28 : _GEN_3565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3567 = 8'hef == io_data_in[103:96] ? 8'hdf : _GEN_3566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3568 = 8'hf0 == io_data_in[103:96] ? 8'h8c : _GEN_3567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3569 = 8'hf1 == io_data_in[103:96] ? 8'ha1 : _GEN_3568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3570 = 8'hf2 == io_data_in[103:96] ? 8'h89 : _GEN_3569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3571 = 8'hf3 == io_data_in[103:96] ? 8'hd : _GEN_3570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3572 = 8'hf4 == io_data_in[103:96] ? 8'hbf : _GEN_3571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3573 = 8'hf5 == io_data_in[103:96] ? 8'he6 : _GEN_3572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3574 = 8'hf6 == io_data_in[103:96] ? 8'h42 : _GEN_3573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3575 = 8'hf7 == io_data_in[103:96] ? 8'h68 : _GEN_3574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3576 = 8'hf8 == io_data_in[103:96] ? 8'h41 : _GEN_3575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3577 = 8'hf9 == io_data_in[103:96] ? 8'h99 : _GEN_3576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3578 = 8'hfa == io_data_in[103:96] ? 8'h2d : _GEN_3577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3579 = 8'hfb == io_data_in[103:96] ? 8'hf : _GEN_3578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3580 = 8'hfc == io_data_in[103:96] ? 8'hb0 : _GEN_3579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3581 = 8'hfd == io_data_in[103:96] ? 8'h54 : _GEN_3580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3582 = 8'hfe == io_data_in[103:96] ? 8'hbb : _GEN_3581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3583 = 8'hff == io_data_in[103:96] ? 8'h16 : _GEN_3582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3585 = 8'h1 == io_data_in[127:120] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3586 = 8'h2 == io_data_in[127:120] ? 8'h77 : _GEN_3585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3587 = 8'h3 == io_data_in[127:120] ? 8'h7b : _GEN_3586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3588 = 8'h4 == io_data_in[127:120] ? 8'hf2 : _GEN_3587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3589 = 8'h5 == io_data_in[127:120] ? 8'h6b : _GEN_3588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3590 = 8'h6 == io_data_in[127:120] ? 8'h6f : _GEN_3589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3591 = 8'h7 == io_data_in[127:120] ? 8'hc5 : _GEN_3590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3592 = 8'h8 == io_data_in[127:120] ? 8'h30 : _GEN_3591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3593 = 8'h9 == io_data_in[127:120] ? 8'h1 : _GEN_3592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3594 = 8'ha == io_data_in[127:120] ? 8'h67 : _GEN_3593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3595 = 8'hb == io_data_in[127:120] ? 8'h2b : _GEN_3594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3596 = 8'hc == io_data_in[127:120] ? 8'hfe : _GEN_3595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3597 = 8'hd == io_data_in[127:120] ? 8'hd7 : _GEN_3596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3598 = 8'he == io_data_in[127:120] ? 8'hab : _GEN_3597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3599 = 8'hf == io_data_in[127:120] ? 8'h76 : _GEN_3598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3600 = 8'h10 == io_data_in[127:120] ? 8'hca : _GEN_3599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3601 = 8'h11 == io_data_in[127:120] ? 8'h82 : _GEN_3600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3602 = 8'h12 == io_data_in[127:120] ? 8'hc9 : _GEN_3601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3603 = 8'h13 == io_data_in[127:120] ? 8'h7d : _GEN_3602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3604 = 8'h14 == io_data_in[127:120] ? 8'hfa : _GEN_3603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3605 = 8'h15 == io_data_in[127:120] ? 8'h59 : _GEN_3604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3606 = 8'h16 == io_data_in[127:120] ? 8'h47 : _GEN_3605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3607 = 8'h17 == io_data_in[127:120] ? 8'hf0 : _GEN_3606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3608 = 8'h18 == io_data_in[127:120] ? 8'had : _GEN_3607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3609 = 8'h19 == io_data_in[127:120] ? 8'hd4 : _GEN_3608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3610 = 8'h1a == io_data_in[127:120] ? 8'ha2 : _GEN_3609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3611 = 8'h1b == io_data_in[127:120] ? 8'haf : _GEN_3610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3612 = 8'h1c == io_data_in[127:120] ? 8'h9c : _GEN_3611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3613 = 8'h1d == io_data_in[127:120] ? 8'ha4 : _GEN_3612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3614 = 8'h1e == io_data_in[127:120] ? 8'h72 : _GEN_3613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3615 = 8'h1f == io_data_in[127:120] ? 8'hc0 : _GEN_3614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3616 = 8'h20 == io_data_in[127:120] ? 8'hb7 : _GEN_3615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3617 = 8'h21 == io_data_in[127:120] ? 8'hfd : _GEN_3616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3618 = 8'h22 == io_data_in[127:120] ? 8'h93 : _GEN_3617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3619 = 8'h23 == io_data_in[127:120] ? 8'h26 : _GEN_3618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3620 = 8'h24 == io_data_in[127:120] ? 8'h36 : _GEN_3619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3621 = 8'h25 == io_data_in[127:120] ? 8'h3f : _GEN_3620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3622 = 8'h26 == io_data_in[127:120] ? 8'hf7 : _GEN_3621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3623 = 8'h27 == io_data_in[127:120] ? 8'hcc : _GEN_3622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3624 = 8'h28 == io_data_in[127:120] ? 8'h34 : _GEN_3623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3625 = 8'h29 == io_data_in[127:120] ? 8'ha5 : _GEN_3624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3626 = 8'h2a == io_data_in[127:120] ? 8'he5 : _GEN_3625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3627 = 8'h2b == io_data_in[127:120] ? 8'hf1 : _GEN_3626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3628 = 8'h2c == io_data_in[127:120] ? 8'h71 : _GEN_3627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3629 = 8'h2d == io_data_in[127:120] ? 8'hd8 : _GEN_3628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3630 = 8'h2e == io_data_in[127:120] ? 8'h31 : _GEN_3629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3631 = 8'h2f == io_data_in[127:120] ? 8'h15 : _GEN_3630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3632 = 8'h30 == io_data_in[127:120] ? 8'h4 : _GEN_3631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3633 = 8'h31 == io_data_in[127:120] ? 8'hc7 : _GEN_3632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3634 = 8'h32 == io_data_in[127:120] ? 8'h23 : _GEN_3633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3635 = 8'h33 == io_data_in[127:120] ? 8'hc3 : _GEN_3634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3636 = 8'h34 == io_data_in[127:120] ? 8'h18 : _GEN_3635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3637 = 8'h35 == io_data_in[127:120] ? 8'h96 : _GEN_3636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3638 = 8'h36 == io_data_in[127:120] ? 8'h5 : _GEN_3637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3639 = 8'h37 == io_data_in[127:120] ? 8'h9a : _GEN_3638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3640 = 8'h38 == io_data_in[127:120] ? 8'h7 : _GEN_3639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3641 = 8'h39 == io_data_in[127:120] ? 8'h12 : _GEN_3640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3642 = 8'h3a == io_data_in[127:120] ? 8'h80 : _GEN_3641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3643 = 8'h3b == io_data_in[127:120] ? 8'he2 : _GEN_3642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3644 = 8'h3c == io_data_in[127:120] ? 8'heb : _GEN_3643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3645 = 8'h3d == io_data_in[127:120] ? 8'h27 : _GEN_3644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3646 = 8'h3e == io_data_in[127:120] ? 8'hb2 : _GEN_3645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3647 = 8'h3f == io_data_in[127:120] ? 8'h75 : _GEN_3646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3648 = 8'h40 == io_data_in[127:120] ? 8'h9 : _GEN_3647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3649 = 8'h41 == io_data_in[127:120] ? 8'h83 : _GEN_3648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3650 = 8'h42 == io_data_in[127:120] ? 8'h2c : _GEN_3649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3651 = 8'h43 == io_data_in[127:120] ? 8'h1a : _GEN_3650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3652 = 8'h44 == io_data_in[127:120] ? 8'h1b : _GEN_3651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3653 = 8'h45 == io_data_in[127:120] ? 8'h6e : _GEN_3652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3654 = 8'h46 == io_data_in[127:120] ? 8'h5a : _GEN_3653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3655 = 8'h47 == io_data_in[127:120] ? 8'ha0 : _GEN_3654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3656 = 8'h48 == io_data_in[127:120] ? 8'h52 : _GEN_3655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3657 = 8'h49 == io_data_in[127:120] ? 8'h3b : _GEN_3656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3658 = 8'h4a == io_data_in[127:120] ? 8'hd6 : _GEN_3657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3659 = 8'h4b == io_data_in[127:120] ? 8'hb3 : _GEN_3658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3660 = 8'h4c == io_data_in[127:120] ? 8'h29 : _GEN_3659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3661 = 8'h4d == io_data_in[127:120] ? 8'he3 : _GEN_3660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3662 = 8'h4e == io_data_in[127:120] ? 8'h2f : _GEN_3661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3663 = 8'h4f == io_data_in[127:120] ? 8'h84 : _GEN_3662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3664 = 8'h50 == io_data_in[127:120] ? 8'h53 : _GEN_3663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3665 = 8'h51 == io_data_in[127:120] ? 8'hd1 : _GEN_3664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3666 = 8'h52 == io_data_in[127:120] ? 8'h0 : _GEN_3665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3667 = 8'h53 == io_data_in[127:120] ? 8'hed : _GEN_3666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3668 = 8'h54 == io_data_in[127:120] ? 8'h20 : _GEN_3667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3669 = 8'h55 == io_data_in[127:120] ? 8'hfc : _GEN_3668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3670 = 8'h56 == io_data_in[127:120] ? 8'hb1 : _GEN_3669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3671 = 8'h57 == io_data_in[127:120] ? 8'h5b : _GEN_3670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3672 = 8'h58 == io_data_in[127:120] ? 8'h6a : _GEN_3671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3673 = 8'h59 == io_data_in[127:120] ? 8'hcb : _GEN_3672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3674 = 8'h5a == io_data_in[127:120] ? 8'hbe : _GEN_3673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3675 = 8'h5b == io_data_in[127:120] ? 8'h39 : _GEN_3674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3676 = 8'h5c == io_data_in[127:120] ? 8'h4a : _GEN_3675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3677 = 8'h5d == io_data_in[127:120] ? 8'h4c : _GEN_3676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3678 = 8'h5e == io_data_in[127:120] ? 8'h58 : _GEN_3677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3679 = 8'h5f == io_data_in[127:120] ? 8'hcf : _GEN_3678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3680 = 8'h60 == io_data_in[127:120] ? 8'hd0 : _GEN_3679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3681 = 8'h61 == io_data_in[127:120] ? 8'hef : _GEN_3680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3682 = 8'h62 == io_data_in[127:120] ? 8'haa : _GEN_3681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3683 = 8'h63 == io_data_in[127:120] ? 8'hfb : _GEN_3682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3684 = 8'h64 == io_data_in[127:120] ? 8'h43 : _GEN_3683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3685 = 8'h65 == io_data_in[127:120] ? 8'h4d : _GEN_3684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3686 = 8'h66 == io_data_in[127:120] ? 8'h33 : _GEN_3685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3687 = 8'h67 == io_data_in[127:120] ? 8'h85 : _GEN_3686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3688 = 8'h68 == io_data_in[127:120] ? 8'h45 : _GEN_3687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3689 = 8'h69 == io_data_in[127:120] ? 8'hf9 : _GEN_3688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3690 = 8'h6a == io_data_in[127:120] ? 8'h2 : _GEN_3689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3691 = 8'h6b == io_data_in[127:120] ? 8'h7f : _GEN_3690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3692 = 8'h6c == io_data_in[127:120] ? 8'h50 : _GEN_3691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3693 = 8'h6d == io_data_in[127:120] ? 8'h3c : _GEN_3692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3694 = 8'h6e == io_data_in[127:120] ? 8'h9f : _GEN_3693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3695 = 8'h6f == io_data_in[127:120] ? 8'ha8 : _GEN_3694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3696 = 8'h70 == io_data_in[127:120] ? 8'h51 : _GEN_3695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3697 = 8'h71 == io_data_in[127:120] ? 8'ha3 : _GEN_3696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3698 = 8'h72 == io_data_in[127:120] ? 8'h40 : _GEN_3697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3699 = 8'h73 == io_data_in[127:120] ? 8'h8f : _GEN_3698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3700 = 8'h74 == io_data_in[127:120] ? 8'h92 : _GEN_3699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3701 = 8'h75 == io_data_in[127:120] ? 8'h9d : _GEN_3700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3702 = 8'h76 == io_data_in[127:120] ? 8'h38 : _GEN_3701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3703 = 8'h77 == io_data_in[127:120] ? 8'hf5 : _GEN_3702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3704 = 8'h78 == io_data_in[127:120] ? 8'hbc : _GEN_3703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3705 = 8'h79 == io_data_in[127:120] ? 8'hb6 : _GEN_3704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3706 = 8'h7a == io_data_in[127:120] ? 8'hda : _GEN_3705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3707 = 8'h7b == io_data_in[127:120] ? 8'h21 : _GEN_3706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3708 = 8'h7c == io_data_in[127:120] ? 8'h10 : _GEN_3707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3709 = 8'h7d == io_data_in[127:120] ? 8'hff : _GEN_3708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3710 = 8'h7e == io_data_in[127:120] ? 8'hf3 : _GEN_3709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3711 = 8'h7f == io_data_in[127:120] ? 8'hd2 : _GEN_3710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3712 = 8'h80 == io_data_in[127:120] ? 8'hcd : _GEN_3711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3713 = 8'h81 == io_data_in[127:120] ? 8'hc : _GEN_3712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3714 = 8'h82 == io_data_in[127:120] ? 8'h13 : _GEN_3713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3715 = 8'h83 == io_data_in[127:120] ? 8'hec : _GEN_3714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3716 = 8'h84 == io_data_in[127:120] ? 8'h5f : _GEN_3715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3717 = 8'h85 == io_data_in[127:120] ? 8'h97 : _GEN_3716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3718 = 8'h86 == io_data_in[127:120] ? 8'h44 : _GEN_3717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3719 = 8'h87 == io_data_in[127:120] ? 8'h17 : _GEN_3718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3720 = 8'h88 == io_data_in[127:120] ? 8'hc4 : _GEN_3719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3721 = 8'h89 == io_data_in[127:120] ? 8'ha7 : _GEN_3720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3722 = 8'h8a == io_data_in[127:120] ? 8'h7e : _GEN_3721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3723 = 8'h8b == io_data_in[127:120] ? 8'h3d : _GEN_3722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3724 = 8'h8c == io_data_in[127:120] ? 8'h64 : _GEN_3723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3725 = 8'h8d == io_data_in[127:120] ? 8'h5d : _GEN_3724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3726 = 8'h8e == io_data_in[127:120] ? 8'h19 : _GEN_3725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3727 = 8'h8f == io_data_in[127:120] ? 8'h73 : _GEN_3726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3728 = 8'h90 == io_data_in[127:120] ? 8'h60 : _GEN_3727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3729 = 8'h91 == io_data_in[127:120] ? 8'h81 : _GEN_3728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3730 = 8'h92 == io_data_in[127:120] ? 8'h4f : _GEN_3729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3731 = 8'h93 == io_data_in[127:120] ? 8'hdc : _GEN_3730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3732 = 8'h94 == io_data_in[127:120] ? 8'h22 : _GEN_3731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3733 = 8'h95 == io_data_in[127:120] ? 8'h2a : _GEN_3732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3734 = 8'h96 == io_data_in[127:120] ? 8'h90 : _GEN_3733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3735 = 8'h97 == io_data_in[127:120] ? 8'h88 : _GEN_3734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3736 = 8'h98 == io_data_in[127:120] ? 8'h46 : _GEN_3735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3737 = 8'h99 == io_data_in[127:120] ? 8'hee : _GEN_3736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3738 = 8'h9a == io_data_in[127:120] ? 8'hb8 : _GEN_3737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3739 = 8'h9b == io_data_in[127:120] ? 8'h14 : _GEN_3738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3740 = 8'h9c == io_data_in[127:120] ? 8'hde : _GEN_3739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3741 = 8'h9d == io_data_in[127:120] ? 8'h5e : _GEN_3740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3742 = 8'h9e == io_data_in[127:120] ? 8'hb : _GEN_3741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3743 = 8'h9f == io_data_in[127:120] ? 8'hdb : _GEN_3742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3744 = 8'ha0 == io_data_in[127:120] ? 8'he0 : _GEN_3743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3745 = 8'ha1 == io_data_in[127:120] ? 8'h32 : _GEN_3744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3746 = 8'ha2 == io_data_in[127:120] ? 8'h3a : _GEN_3745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3747 = 8'ha3 == io_data_in[127:120] ? 8'ha : _GEN_3746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3748 = 8'ha4 == io_data_in[127:120] ? 8'h49 : _GEN_3747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3749 = 8'ha5 == io_data_in[127:120] ? 8'h6 : _GEN_3748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3750 = 8'ha6 == io_data_in[127:120] ? 8'h24 : _GEN_3749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3751 = 8'ha7 == io_data_in[127:120] ? 8'h5c : _GEN_3750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3752 = 8'ha8 == io_data_in[127:120] ? 8'hc2 : _GEN_3751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3753 = 8'ha9 == io_data_in[127:120] ? 8'hd3 : _GEN_3752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3754 = 8'haa == io_data_in[127:120] ? 8'hac : _GEN_3753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3755 = 8'hab == io_data_in[127:120] ? 8'h62 : _GEN_3754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3756 = 8'hac == io_data_in[127:120] ? 8'h91 : _GEN_3755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3757 = 8'had == io_data_in[127:120] ? 8'h95 : _GEN_3756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3758 = 8'hae == io_data_in[127:120] ? 8'he4 : _GEN_3757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3759 = 8'haf == io_data_in[127:120] ? 8'h79 : _GEN_3758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3760 = 8'hb0 == io_data_in[127:120] ? 8'he7 : _GEN_3759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3761 = 8'hb1 == io_data_in[127:120] ? 8'hc8 : _GEN_3760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3762 = 8'hb2 == io_data_in[127:120] ? 8'h37 : _GEN_3761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3763 = 8'hb3 == io_data_in[127:120] ? 8'h6d : _GEN_3762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3764 = 8'hb4 == io_data_in[127:120] ? 8'h8d : _GEN_3763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3765 = 8'hb5 == io_data_in[127:120] ? 8'hd5 : _GEN_3764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3766 = 8'hb6 == io_data_in[127:120] ? 8'h4e : _GEN_3765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3767 = 8'hb7 == io_data_in[127:120] ? 8'ha9 : _GEN_3766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3768 = 8'hb8 == io_data_in[127:120] ? 8'h6c : _GEN_3767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3769 = 8'hb9 == io_data_in[127:120] ? 8'h56 : _GEN_3768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3770 = 8'hba == io_data_in[127:120] ? 8'hf4 : _GEN_3769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3771 = 8'hbb == io_data_in[127:120] ? 8'hea : _GEN_3770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3772 = 8'hbc == io_data_in[127:120] ? 8'h65 : _GEN_3771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3773 = 8'hbd == io_data_in[127:120] ? 8'h7a : _GEN_3772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3774 = 8'hbe == io_data_in[127:120] ? 8'hae : _GEN_3773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3775 = 8'hbf == io_data_in[127:120] ? 8'h8 : _GEN_3774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3776 = 8'hc0 == io_data_in[127:120] ? 8'hba : _GEN_3775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3777 = 8'hc1 == io_data_in[127:120] ? 8'h78 : _GEN_3776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3778 = 8'hc2 == io_data_in[127:120] ? 8'h25 : _GEN_3777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3779 = 8'hc3 == io_data_in[127:120] ? 8'h2e : _GEN_3778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3780 = 8'hc4 == io_data_in[127:120] ? 8'h1c : _GEN_3779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3781 = 8'hc5 == io_data_in[127:120] ? 8'ha6 : _GEN_3780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3782 = 8'hc6 == io_data_in[127:120] ? 8'hb4 : _GEN_3781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3783 = 8'hc7 == io_data_in[127:120] ? 8'hc6 : _GEN_3782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3784 = 8'hc8 == io_data_in[127:120] ? 8'he8 : _GEN_3783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3785 = 8'hc9 == io_data_in[127:120] ? 8'hdd : _GEN_3784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3786 = 8'hca == io_data_in[127:120] ? 8'h74 : _GEN_3785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3787 = 8'hcb == io_data_in[127:120] ? 8'h1f : _GEN_3786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3788 = 8'hcc == io_data_in[127:120] ? 8'h4b : _GEN_3787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3789 = 8'hcd == io_data_in[127:120] ? 8'hbd : _GEN_3788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3790 = 8'hce == io_data_in[127:120] ? 8'h8b : _GEN_3789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3791 = 8'hcf == io_data_in[127:120] ? 8'h8a : _GEN_3790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3792 = 8'hd0 == io_data_in[127:120] ? 8'h70 : _GEN_3791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3793 = 8'hd1 == io_data_in[127:120] ? 8'h3e : _GEN_3792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3794 = 8'hd2 == io_data_in[127:120] ? 8'hb5 : _GEN_3793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3795 = 8'hd3 == io_data_in[127:120] ? 8'h66 : _GEN_3794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3796 = 8'hd4 == io_data_in[127:120] ? 8'h48 : _GEN_3795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3797 = 8'hd5 == io_data_in[127:120] ? 8'h3 : _GEN_3796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3798 = 8'hd6 == io_data_in[127:120] ? 8'hf6 : _GEN_3797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3799 = 8'hd7 == io_data_in[127:120] ? 8'he : _GEN_3798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3800 = 8'hd8 == io_data_in[127:120] ? 8'h61 : _GEN_3799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3801 = 8'hd9 == io_data_in[127:120] ? 8'h35 : _GEN_3800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3802 = 8'hda == io_data_in[127:120] ? 8'h57 : _GEN_3801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3803 = 8'hdb == io_data_in[127:120] ? 8'hb9 : _GEN_3802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3804 = 8'hdc == io_data_in[127:120] ? 8'h86 : _GEN_3803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3805 = 8'hdd == io_data_in[127:120] ? 8'hc1 : _GEN_3804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3806 = 8'hde == io_data_in[127:120] ? 8'h1d : _GEN_3805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3807 = 8'hdf == io_data_in[127:120] ? 8'h9e : _GEN_3806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3808 = 8'he0 == io_data_in[127:120] ? 8'he1 : _GEN_3807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3809 = 8'he1 == io_data_in[127:120] ? 8'hf8 : _GEN_3808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3810 = 8'he2 == io_data_in[127:120] ? 8'h98 : _GEN_3809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3811 = 8'he3 == io_data_in[127:120] ? 8'h11 : _GEN_3810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3812 = 8'he4 == io_data_in[127:120] ? 8'h69 : _GEN_3811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3813 = 8'he5 == io_data_in[127:120] ? 8'hd9 : _GEN_3812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3814 = 8'he6 == io_data_in[127:120] ? 8'h8e : _GEN_3813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3815 = 8'he7 == io_data_in[127:120] ? 8'h94 : _GEN_3814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3816 = 8'he8 == io_data_in[127:120] ? 8'h9b : _GEN_3815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3817 = 8'he9 == io_data_in[127:120] ? 8'h1e : _GEN_3816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3818 = 8'hea == io_data_in[127:120] ? 8'h87 : _GEN_3817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3819 = 8'heb == io_data_in[127:120] ? 8'he9 : _GEN_3818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3820 = 8'hec == io_data_in[127:120] ? 8'hce : _GEN_3819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3821 = 8'hed == io_data_in[127:120] ? 8'h55 : _GEN_3820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3822 = 8'hee == io_data_in[127:120] ? 8'h28 : _GEN_3821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3823 = 8'hef == io_data_in[127:120] ? 8'hdf : _GEN_3822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3824 = 8'hf0 == io_data_in[127:120] ? 8'h8c : _GEN_3823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3825 = 8'hf1 == io_data_in[127:120] ? 8'ha1 : _GEN_3824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3826 = 8'hf2 == io_data_in[127:120] ? 8'h89 : _GEN_3825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3827 = 8'hf3 == io_data_in[127:120] ? 8'hd : _GEN_3826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3828 = 8'hf4 == io_data_in[127:120] ? 8'hbf : _GEN_3827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3829 = 8'hf5 == io_data_in[127:120] ? 8'he6 : _GEN_3828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3830 = 8'hf6 == io_data_in[127:120] ? 8'h42 : _GEN_3829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3831 = 8'hf7 == io_data_in[127:120] ? 8'h68 : _GEN_3830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3832 = 8'hf8 == io_data_in[127:120] ? 8'h41 : _GEN_3831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3833 = 8'hf9 == io_data_in[127:120] ? 8'h99 : _GEN_3832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3834 = 8'hfa == io_data_in[127:120] ? 8'h2d : _GEN_3833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3835 = 8'hfb == io_data_in[127:120] ? 8'hf : _GEN_3834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3836 = 8'hfc == io_data_in[127:120] ? 8'hb0 : _GEN_3835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3837 = 8'hfd == io_data_in[127:120] ? 8'h54 : _GEN_3836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3838 = 8'hfe == io_data_in[127:120] ? 8'hbb : _GEN_3837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3839 = 8'hff == io_data_in[127:120] ? 8'h16 : _GEN_3838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3841 = 8'h1 == io_data_in[119:112] ? 8'h7c : 8'h63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3842 = 8'h2 == io_data_in[119:112] ? 8'h77 : _GEN_3841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3843 = 8'h3 == io_data_in[119:112] ? 8'h7b : _GEN_3842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3844 = 8'h4 == io_data_in[119:112] ? 8'hf2 : _GEN_3843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3845 = 8'h5 == io_data_in[119:112] ? 8'h6b : _GEN_3844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3846 = 8'h6 == io_data_in[119:112] ? 8'h6f : _GEN_3845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3847 = 8'h7 == io_data_in[119:112] ? 8'hc5 : _GEN_3846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3848 = 8'h8 == io_data_in[119:112] ? 8'h30 : _GEN_3847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3849 = 8'h9 == io_data_in[119:112] ? 8'h1 : _GEN_3848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3850 = 8'ha == io_data_in[119:112] ? 8'h67 : _GEN_3849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3851 = 8'hb == io_data_in[119:112] ? 8'h2b : _GEN_3850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3852 = 8'hc == io_data_in[119:112] ? 8'hfe : _GEN_3851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3853 = 8'hd == io_data_in[119:112] ? 8'hd7 : _GEN_3852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3854 = 8'he == io_data_in[119:112] ? 8'hab : _GEN_3853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3855 = 8'hf == io_data_in[119:112] ? 8'h76 : _GEN_3854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3856 = 8'h10 == io_data_in[119:112] ? 8'hca : _GEN_3855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3857 = 8'h11 == io_data_in[119:112] ? 8'h82 : _GEN_3856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3858 = 8'h12 == io_data_in[119:112] ? 8'hc9 : _GEN_3857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3859 = 8'h13 == io_data_in[119:112] ? 8'h7d : _GEN_3858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3860 = 8'h14 == io_data_in[119:112] ? 8'hfa : _GEN_3859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3861 = 8'h15 == io_data_in[119:112] ? 8'h59 : _GEN_3860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3862 = 8'h16 == io_data_in[119:112] ? 8'h47 : _GEN_3861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3863 = 8'h17 == io_data_in[119:112] ? 8'hf0 : _GEN_3862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3864 = 8'h18 == io_data_in[119:112] ? 8'had : _GEN_3863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3865 = 8'h19 == io_data_in[119:112] ? 8'hd4 : _GEN_3864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3866 = 8'h1a == io_data_in[119:112] ? 8'ha2 : _GEN_3865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3867 = 8'h1b == io_data_in[119:112] ? 8'haf : _GEN_3866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3868 = 8'h1c == io_data_in[119:112] ? 8'h9c : _GEN_3867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3869 = 8'h1d == io_data_in[119:112] ? 8'ha4 : _GEN_3868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3870 = 8'h1e == io_data_in[119:112] ? 8'h72 : _GEN_3869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3871 = 8'h1f == io_data_in[119:112] ? 8'hc0 : _GEN_3870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3872 = 8'h20 == io_data_in[119:112] ? 8'hb7 : _GEN_3871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3873 = 8'h21 == io_data_in[119:112] ? 8'hfd : _GEN_3872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3874 = 8'h22 == io_data_in[119:112] ? 8'h93 : _GEN_3873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3875 = 8'h23 == io_data_in[119:112] ? 8'h26 : _GEN_3874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3876 = 8'h24 == io_data_in[119:112] ? 8'h36 : _GEN_3875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3877 = 8'h25 == io_data_in[119:112] ? 8'h3f : _GEN_3876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3878 = 8'h26 == io_data_in[119:112] ? 8'hf7 : _GEN_3877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3879 = 8'h27 == io_data_in[119:112] ? 8'hcc : _GEN_3878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3880 = 8'h28 == io_data_in[119:112] ? 8'h34 : _GEN_3879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3881 = 8'h29 == io_data_in[119:112] ? 8'ha5 : _GEN_3880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3882 = 8'h2a == io_data_in[119:112] ? 8'he5 : _GEN_3881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3883 = 8'h2b == io_data_in[119:112] ? 8'hf1 : _GEN_3882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3884 = 8'h2c == io_data_in[119:112] ? 8'h71 : _GEN_3883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3885 = 8'h2d == io_data_in[119:112] ? 8'hd8 : _GEN_3884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3886 = 8'h2e == io_data_in[119:112] ? 8'h31 : _GEN_3885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3887 = 8'h2f == io_data_in[119:112] ? 8'h15 : _GEN_3886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3888 = 8'h30 == io_data_in[119:112] ? 8'h4 : _GEN_3887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3889 = 8'h31 == io_data_in[119:112] ? 8'hc7 : _GEN_3888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3890 = 8'h32 == io_data_in[119:112] ? 8'h23 : _GEN_3889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3891 = 8'h33 == io_data_in[119:112] ? 8'hc3 : _GEN_3890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3892 = 8'h34 == io_data_in[119:112] ? 8'h18 : _GEN_3891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3893 = 8'h35 == io_data_in[119:112] ? 8'h96 : _GEN_3892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3894 = 8'h36 == io_data_in[119:112] ? 8'h5 : _GEN_3893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3895 = 8'h37 == io_data_in[119:112] ? 8'h9a : _GEN_3894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3896 = 8'h38 == io_data_in[119:112] ? 8'h7 : _GEN_3895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3897 = 8'h39 == io_data_in[119:112] ? 8'h12 : _GEN_3896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3898 = 8'h3a == io_data_in[119:112] ? 8'h80 : _GEN_3897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3899 = 8'h3b == io_data_in[119:112] ? 8'he2 : _GEN_3898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3900 = 8'h3c == io_data_in[119:112] ? 8'heb : _GEN_3899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3901 = 8'h3d == io_data_in[119:112] ? 8'h27 : _GEN_3900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3902 = 8'h3e == io_data_in[119:112] ? 8'hb2 : _GEN_3901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3903 = 8'h3f == io_data_in[119:112] ? 8'h75 : _GEN_3902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3904 = 8'h40 == io_data_in[119:112] ? 8'h9 : _GEN_3903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3905 = 8'h41 == io_data_in[119:112] ? 8'h83 : _GEN_3904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3906 = 8'h42 == io_data_in[119:112] ? 8'h2c : _GEN_3905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3907 = 8'h43 == io_data_in[119:112] ? 8'h1a : _GEN_3906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3908 = 8'h44 == io_data_in[119:112] ? 8'h1b : _GEN_3907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3909 = 8'h45 == io_data_in[119:112] ? 8'h6e : _GEN_3908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3910 = 8'h46 == io_data_in[119:112] ? 8'h5a : _GEN_3909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3911 = 8'h47 == io_data_in[119:112] ? 8'ha0 : _GEN_3910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3912 = 8'h48 == io_data_in[119:112] ? 8'h52 : _GEN_3911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3913 = 8'h49 == io_data_in[119:112] ? 8'h3b : _GEN_3912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3914 = 8'h4a == io_data_in[119:112] ? 8'hd6 : _GEN_3913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3915 = 8'h4b == io_data_in[119:112] ? 8'hb3 : _GEN_3914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3916 = 8'h4c == io_data_in[119:112] ? 8'h29 : _GEN_3915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3917 = 8'h4d == io_data_in[119:112] ? 8'he3 : _GEN_3916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3918 = 8'h4e == io_data_in[119:112] ? 8'h2f : _GEN_3917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3919 = 8'h4f == io_data_in[119:112] ? 8'h84 : _GEN_3918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3920 = 8'h50 == io_data_in[119:112] ? 8'h53 : _GEN_3919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3921 = 8'h51 == io_data_in[119:112] ? 8'hd1 : _GEN_3920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3922 = 8'h52 == io_data_in[119:112] ? 8'h0 : _GEN_3921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3923 = 8'h53 == io_data_in[119:112] ? 8'hed : _GEN_3922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3924 = 8'h54 == io_data_in[119:112] ? 8'h20 : _GEN_3923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3925 = 8'h55 == io_data_in[119:112] ? 8'hfc : _GEN_3924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3926 = 8'h56 == io_data_in[119:112] ? 8'hb1 : _GEN_3925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3927 = 8'h57 == io_data_in[119:112] ? 8'h5b : _GEN_3926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3928 = 8'h58 == io_data_in[119:112] ? 8'h6a : _GEN_3927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3929 = 8'h59 == io_data_in[119:112] ? 8'hcb : _GEN_3928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3930 = 8'h5a == io_data_in[119:112] ? 8'hbe : _GEN_3929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3931 = 8'h5b == io_data_in[119:112] ? 8'h39 : _GEN_3930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3932 = 8'h5c == io_data_in[119:112] ? 8'h4a : _GEN_3931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3933 = 8'h5d == io_data_in[119:112] ? 8'h4c : _GEN_3932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3934 = 8'h5e == io_data_in[119:112] ? 8'h58 : _GEN_3933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3935 = 8'h5f == io_data_in[119:112] ? 8'hcf : _GEN_3934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3936 = 8'h60 == io_data_in[119:112] ? 8'hd0 : _GEN_3935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3937 = 8'h61 == io_data_in[119:112] ? 8'hef : _GEN_3936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3938 = 8'h62 == io_data_in[119:112] ? 8'haa : _GEN_3937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3939 = 8'h63 == io_data_in[119:112] ? 8'hfb : _GEN_3938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3940 = 8'h64 == io_data_in[119:112] ? 8'h43 : _GEN_3939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3941 = 8'h65 == io_data_in[119:112] ? 8'h4d : _GEN_3940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3942 = 8'h66 == io_data_in[119:112] ? 8'h33 : _GEN_3941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3943 = 8'h67 == io_data_in[119:112] ? 8'h85 : _GEN_3942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3944 = 8'h68 == io_data_in[119:112] ? 8'h45 : _GEN_3943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3945 = 8'h69 == io_data_in[119:112] ? 8'hf9 : _GEN_3944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3946 = 8'h6a == io_data_in[119:112] ? 8'h2 : _GEN_3945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3947 = 8'h6b == io_data_in[119:112] ? 8'h7f : _GEN_3946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3948 = 8'h6c == io_data_in[119:112] ? 8'h50 : _GEN_3947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3949 = 8'h6d == io_data_in[119:112] ? 8'h3c : _GEN_3948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3950 = 8'h6e == io_data_in[119:112] ? 8'h9f : _GEN_3949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3951 = 8'h6f == io_data_in[119:112] ? 8'ha8 : _GEN_3950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3952 = 8'h70 == io_data_in[119:112] ? 8'h51 : _GEN_3951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3953 = 8'h71 == io_data_in[119:112] ? 8'ha3 : _GEN_3952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3954 = 8'h72 == io_data_in[119:112] ? 8'h40 : _GEN_3953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3955 = 8'h73 == io_data_in[119:112] ? 8'h8f : _GEN_3954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3956 = 8'h74 == io_data_in[119:112] ? 8'h92 : _GEN_3955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3957 = 8'h75 == io_data_in[119:112] ? 8'h9d : _GEN_3956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3958 = 8'h76 == io_data_in[119:112] ? 8'h38 : _GEN_3957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3959 = 8'h77 == io_data_in[119:112] ? 8'hf5 : _GEN_3958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3960 = 8'h78 == io_data_in[119:112] ? 8'hbc : _GEN_3959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3961 = 8'h79 == io_data_in[119:112] ? 8'hb6 : _GEN_3960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3962 = 8'h7a == io_data_in[119:112] ? 8'hda : _GEN_3961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3963 = 8'h7b == io_data_in[119:112] ? 8'h21 : _GEN_3962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3964 = 8'h7c == io_data_in[119:112] ? 8'h10 : _GEN_3963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3965 = 8'h7d == io_data_in[119:112] ? 8'hff : _GEN_3964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3966 = 8'h7e == io_data_in[119:112] ? 8'hf3 : _GEN_3965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3967 = 8'h7f == io_data_in[119:112] ? 8'hd2 : _GEN_3966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3968 = 8'h80 == io_data_in[119:112] ? 8'hcd : _GEN_3967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3969 = 8'h81 == io_data_in[119:112] ? 8'hc : _GEN_3968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3970 = 8'h82 == io_data_in[119:112] ? 8'h13 : _GEN_3969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3971 = 8'h83 == io_data_in[119:112] ? 8'hec : _GEN_3970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3972 = 8'h84 == io_data_in[119:112] ? 8'h5f : _GEN_3971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3973 = 8'h85 == io_data_in[119:112] ? 8'h97 : _GEN_3972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3974 = 8'h86 == io_data_in[119:112] ? 8'h44 : _GEN_3973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3975 = 8'h87 == io_data_in[119:112] ? 8'h17 : _GEN_3974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3976 = 8'h88 == io_data_in[119:112] ? 8'hc4 : _GEN_3975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3977 = 8'h89 == io_data_in[119:112] ? 8'ha7 : _GEN_3976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3978 = 8'h8a == io_data_in[119:112] ? 8'h7e : _GEN_3977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3979 = 8'h8b == io_data_in[119:112] ? 8'h3d : _GEN_3978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3980 = 8'h8c == io_data_in[119:112] ? 8'h64 : _GEN_3979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3981 = 8'h8d == io_data_in[119:112] ? 8'h5d : _GEN_3980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3982 = 8'h8e == io_data_in[119:112] ? 8'h19 : _GEN_3981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3983 = 8'h8f == io_data_in[119:112] ? 8'h73 : _GEN_3982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3984 = 8'h90 == io_data_in[119:112] ? 8'h60 : _GEN_3983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3985 = 8'h91 == io_data_in[119:112] ? 8'h81 : _GEN_3984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3986 = 8'h92 == io_data_in[119:112] ? 8'h4f : _GEN_3985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3987 = 8'h93 == io_data_in[119:112] ? 8'hdc : _GEN_3986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3988 = 8'h94 == io_data_in[119:112] ? 8'h22 : _GEN_3987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3989 = 8'h95 == io_data_in[119:112] ? 8'h2a : _GEN_3988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3990 = 8'h96 == io_data_in[119:112] ? 8'h90 : _GEN_3989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3991 = 8'h97 == io_data_in[119:112] ? 8'h88 : _GEN_3990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3992 = 8'h98 == io_data_in[119:112] ? 8'h46 : _GEN_3991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3993 = 8'h99 == io_data_in[119:112] ? 8'hee : _GEN_3992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3994 = 8'h9a == io_data_in[119:112] ? 8'hb8 : _GEN_3993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3995 = 8'h9b == io_data_in[119:112] ? 8'h14 : _GEN_3994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3996 = 8'h9c == io_data_in[119:112] ? 8'hde : _GEN_3995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3997 = 8'h9d == io_data_in[119:112] ? 8'h5e : _GEN_3996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3998 = 8'h9e == io_data_in[119:112] ? 8'hb : _GEN_3997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3999 = 8'h9f == io_data_in[119:112] ? 8'hdb : _GEN_3998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4000 = 8'ha0 == io_data_in[119:112] ? 8'he0 : _GEN_3999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4001 = 8'ha1 == io_data_in[119:112] ? 8'h32 : _GEN_4000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4002 = 8'ha2 == io_data_in[119:112] ? 8'h3a : _GEN_4001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4003 = 8'ha3 == io_data_in[119:112] ? 8'ha : _GEN_4002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4004 = 8'ha4 == io_data_in[119:112] ? 8'h49 : _GEN_4003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4005 = 8'ha5 == io_data_in[119:112] ? 8'h6 : _GEN_4004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4006 = 8'ha6 == io_data_in[119:112] ? 8'h24 : _GEN_4005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4007 = 8'ha7 == io_data_in[119:112] ? 8'h5c : _GEN_4006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4008 = 8'ha8 == io_data_in[119:112] ? 8'hc2 : _GEN_4007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4009 = 8'ha9 == io_data_in[119:112] ? 8'hd3 : _GEN_4008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4010 = 8'haa == io_data_in[119:112] ? 8'hac : _GEN_4009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4011 = 8'hab == io_data_in[119:112] ? 8'h62 : _GEN_4010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4012 = 8'hac == io_data_in[119:112] ? 8'h91 : _GEN_4011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4013 = 8'had == io_data_in[119:112] ? 8'h95 : _GEN_4012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4014 = 8'hae == io_data_in[119:112] ? 8'he4 : _GEN_4013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4015 = 8'haf == io_data_in[119:112] ? 8'h79 : _GEN_4014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4016 = 8'hb0 == io_data_in[119:112] ? 8'he7 : _GEN_4015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4017 = 8'hb1 == io_data_in[119:112] ? 8'hc8 : _GEN_4016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4018 = 8'hb2 == io_data_in[119:112] ? 8'h37 : _GEN_4017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4019 = 8'hb3 == io_data_in[119:112] ? 8'h6d : _GEN_4018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4020 = 8'hb4 == io_data_in[119:112] ? 8'h8d : _GEN_4019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4021 = 8'hb5 == io_data_in[119:112] ? 8'hd5 : _GEN_4020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4022 = 8'hb6 == io_data_in[119:112] ? 8'h4e : _GEN_4021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4023 = 8'hb7 == io_data_in[119:112] ? 8'ha9 : _GEN_4022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4024 = 8'hb8 == io_data_in[119:112] ? 8'h6c : _GEN_4023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4025 = 8'hb9 == io_data_in[119:112] ? 8'h56 : _GEN_4024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4026 = 8'hba == io_data_in[119:112] ? 8'hf4 : _GEN_4025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4027 = 8'hbb == io_data_in[119:112] ? 8'hea : _GEN_4026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4028 = 8'hbc == io_data_in[119:112] ? 8'h65 : _GEN_4027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4029 = 8'hbd == io_data_in[119:112] ? 8'h7a : _GEN_4028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4030 = 8'hbe == io_data_in[119:112] ? 8'hae : _GEN_4029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4031 = 8'hbf == io_data_in[119:112] ? 8'h8 : _GEN_4030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4032 = 8'hc0 == io_data_in[119:112] ? 8'hba : _GEN_4031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4033 = 8'hc1 == io_data_in[119:112] ? 8'h78 : _GEN_4032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4034 = 8'hc2 == io_data_in[119:112] ? 8'h25 : _GEN_4033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4035 = 8'hc3 == io_data_in[119:112] ? 8'h2e : _GEN_4034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4036 = 8'hc4 == io_data_in[119:112] ? 8'h1c : _GEN_4035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4037 = 8'hc5 == io_data_in[119:112] ? 8'ha6 : _GEN_4036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4038 = 8'hc6 == io_data_in[119:112] ? 8'hb4 : _GEN_4037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4039 = 8'hc7 == io_data_in[119:112] ? 8'hc6 : _GEN_4038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4040 = 8'hc8 == io_data_in[119:112] ? 8'he8 : _GEN_4039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4041 = 8'hc9 == io_data_in[119:112] ? 8'hdd : _GEN_4040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4042 = 8'hca == io_data_in[119:112] ? 8'h74 : _GEN_4041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4043 = 8'hcb == io_data_in[119:112] ? 8'h1f : _GEN_4042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4044 = 8'hcc == io_data_in[119:112] ? 8'h4b : _GEN_4043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4045 = 8'hcd == io_data_in[119:112] ? 8'hbd : _GEN_4044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4046 = 8'hce == io_data_in[119:112] ? 8'h8b : _GEN_4045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4047 = 8'hcf == io_data_in[119:112] ? 8'h8a : _GEN_4046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4048 = 8'hd0 == io_data_in[119:112] ? 8'h70 : _GEN_4047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4049 = 8'hd1 == io_data_in[119:112] ? 8'h3e : _GEN_4048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4050 = 8'hd2 == io_data_in[119:112] ? 8'hb5 : _GEN_4049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4051 = 8'hd3 == io_data_in[119:112] ? 8'h66 : _GEN_4050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4052 = 8'hd4 == io_data_in[119:112] ? 8'h48 : _GEN_4051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4053 = 8'hd5 == io_data_in[119:112] ? 8'h3 : _GEN_4052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4054 = 8'hd6 == io_data_in[119:112] ? 8'hf6 : _GEN_4053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4055 = 8'hd7 == io_data_in[119:112] ? 8'he : _GEN_4054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4056 = 8'hd8 == io_data_in[119:112] ? 8'h61 : _GEN_4055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4057 = 8'hd9 == io_data_in[119:112] ? 8'h35 : _GEN_4056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4058 = 8'hda == io_data_in[119:112] ? 8'h57 : _GEN_4057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4059 = 8'hdb == io_data_in[119:112] ? 8'hb9 : _GEN_4058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4060 = 8'hdc == io_data_in[119:112] ? 8'h86 : _GEN_4059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4061 = 8'hdd == io_data_in[119:112] ? 8'hc1 : _GEN_4060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4062 = 8'hde == io_data_in[119:112] ? 8'h1d : _GEN_4061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4063 = 8'hdf == io_data_in[119:112] ? 8'h9e : _GEN_4062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4064 = 8'he0 == io_data_in[119:112] ? 8'he1 : _GEN_4063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4065 = 8'he1 == io_data_in[119:112] ? 8'hf8 : _GEN_4064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4066 = 8'he2 == io_data_in[119:112] ? 8'h98 : _GEN_4065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4067 = 8'he3 == io_data_in[119:112] ? 8'h11 : _GEN_4066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4068 = 8'he4 == io_data_in[119:112] ? 8'h69 : _GEN_4067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4069 = 8'he5 == io_data_in[119:112] ? 8'hd9 : _GEN_4068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4070 = 8'he6 == io_data_in[119:112] ? 8'h8e : _GEN_4069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4071 = 8'he7 == io_data_in[119:112] ? 8'h94 : _GEN_4070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4072 = 8'he8 == io_data_in[119:112] ? 8'h9b : _GEN_4071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4073 = 8'he9 == io_data_in[119:112] ? 8'h1e : _GEN_4072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4074 = 8'hea == io_data_in[119:112] ? 8'h87 : _GEN_4073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4075 = 8'heb == io_data_in[119:112] ? 8'he9 : _GEN_4074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4076 = 8'hec == io_data_in[119:112] ? 8'hce : _GEN_4075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4077 = 8'hed == io_data_in[119:112] ? 8'h55 : _GEN_4076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4078 = 8'hee == io_data_in[119:112] ? 8'h28 : _GEN_4077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4079 = 8'hef == io_data_in[119:112] ? 8'hdf : _GEN_4078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4080 = 8'hf0 == io_data_in[119:112] ? 8'h8c : _GEN_4079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4081 = 8'hf1 == io_data_in[119:112] ? 8'ha1 : _GEN_4080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4082 = 8'hf2 == io_data_in[119:112] ? 8'h89 : _GEN_4081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4083 = 8'hf3 == io_data_in[119:112] ? 8'hd : _GEN_4082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4084 = 8'hf4 == io_data_in[119:112] ? 8'hbf : _GEN_4083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4085 = 8'hf5 == io_data_in[119:112] ? 8'he6 : _GEN_4084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4086 = 8'hf6 == io_data_in[119:112] ? 8'h42 : _GEN_4085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4087 = 8'hf7 == io_data_in[119:112] ? 8'h68 : _GEN_4086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4088 = 8'hf8 == io_data_in[119:112] ? 8'h41 : _GEN_4087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4089 = 8'hf9 == io_data_in[119:112] ? 8'h99 : _GEN_4088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4090 = 8'hfa == io_data_in[119:112] ? 8'h2d : _GEN_4089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4091 = 8'hfb == io_data_in[119:112] ? 8'hf : _GEN_4090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4092 = 8'hfc == io_data_in[119:112] ? 8'hb0 : _GEN_4091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4093 = 8'hfd == io_data_in[119:112] ? 8'h54 : _GEN_4092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4094 = 8'hfe == io_data_in[119:112] ? 8'hbb : _GEN_4093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4095 = 8'hff == io_data_in[119:112] ? 8'h16 : _GEN_4094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [63:0] io_data_out_hi = {_GEN_3839,_GEN_4095,_GEN_3327,_GEN_3583,_GEN_2815,_GEN_3071,_GEN_2303,_GEN_2559}; // @[Cat.scala 30:58]
  assign io_data_out = {io_data_out_hi,io_data_out_lo}; // @[Cat.scala 30:58]
endmodule
/*
module GFMult(
  input  [7:0] io_data_in_1,
  input  [7:0] io_data_in_2,
  output [7:0] io_data_out
);
  wire [10:0] _m_T = {3'h0,io_data_in_1}; // @[Cat.scala 30:58]
  wire  m_hi_hi_hi_hi = io_data_in_2[0]; // @[GFMult.scala 9:58]
  wire [4:0] m_lo = {m_hi_hi_hi_hi,m_hi_hi_hi_hi,m_hi_hi_hi_hi,m_hi_hi_hi_hi,m_hi_hi_hi_hi}; // @[Cat.scala 30:58]
  wire [10:0] _m_T_1 = {m_hi_hi_hi_hi,m_hi_hi_hi_hi,m_hi_hi_hi_hi,m_hi_hi_hi_hi,m_hi_hi_hi_hi,m_hi_hi_hi_hi,m_lo}; // @[Cat.scala 30:58]
  wire [10:0] _m_T_2 = _m_T & _m_T_1; // @[GFMult.scala 9:39]
  wire [10:0] _m_T_3 = {2'h0,io_data_in_1,1'h0}; // @[Cat.scala 30:58]
  wire  m_hi_hi_hi_hi_1 = io_data_in_2[1]; // @[GFMult.scala 10:67]
  wire [4:0] m_lo_1 = {m_hi_hi_hi_hi_1,m_hi_hi_hi_hi_1,m_hi_hi_hi_hi_1,m_hi_hi_hi_hi_1,m_hi_hi_hi_hi_1}; // @[Cat.scala 30:58]
  wire [10:0] _m_T_4 = {m_hi_hi_hi_hi_1,m_hi_hi_hi_hi_1,m_hi_hi_hi_hi_1,m_hi_hi_hi_hi_1,m_hi_hi_hi_hi_1,m_hi_hi_hi_hi_1,
    m_lo_1}; // @[Cat.scala 30:58]
  wire [10:0] _m_T_5 = _m_T_3 & _m_T_4; // @[GFMult.scala 10:48]
  wire [10:0] _m_T_6 = _m_T_2 ^ _m_T_5; // @[GFMult.scala 9:225]
  wire [10:0] _m_T_7 = {1'h0,io_data_in_1,2'h0}; // @[Cat.scala 30:58]
  wire  m_hi_hi_hi_hi_2 = io_data_in_2[2]; // @[GFMult.scala 11:67]
  wire [4:0] m_lo_2 = {m_hi_hi_hi_hi_2,m_hi_hi_hi_hi_2,m_hi_hi_hi_hi_2,m_hi_hi_hi_hi_2,m_hi_hi_hi_hi_2}; // @[Cat.scala 30:58]
  wire [10:0] _m_T_8 = {m_hi_hi_hi_hi_2,m_hi_hi_hi_hi_2,m_hi_hi_hi_hi_2,m_hi_hi_hi_hi_2,m_hi_hi_hi_hi_2,m_hi_hi_hi_hi_2,
    m_lo_2}; // @[Cat.scala 30:58]
  wire [10:0] _m_T_9 = _m_T_7 & _m_T_8; // @[GFMult.scala 11:48]
  wire [10:0] _m_T_10 = _m_T_6 ^ _m_T_9; // @[GFMult.scala 10:234]
  wire [10:0] _m_T_11 = {io_data_in_1,3'h0}; // @[Cat.scala 30:58]
  wire  m_hi_hi_hi_hi_3 = io_data_in_2[3]; // @[GFMult.scala 12:58]
  wire [4:0] m_lo_3 = {m_hi_hi_hi_hi_3,m_hi_hi_hi_hi_3,m_hi_hi_hi_hi_3,m_hi_hi_hi_hi_3,m_hi_hi_hi_hi_3}; // @[Cat.scala 30:58]
  wire [10:0] _m_T_12 = {m_hi_hi_hi_hi_3,m_hi_hi_hi_hi_3,m_hi_hi_hi_hi_3,m_hi_hi_hi_hi_3,m_hi_hi_hi_hi_3,m_hi_hi_hi_hi_3
    ,m_lo_3}; // @[Cat.scala 30:58]
  wire [10:0] _m_T_13 = _m_T_11 & _m_T_12; // @[GFMult.scala 12:39]
  wire [10:0] m = _m_T_10 ^ _m_T_13; // @[GFMult.scala 11:234]
  wire  io_data_out_hi_hi_hi = m[8]; // @[GFMult.scala 13:50]
  wire [7:0] _io_data_out_T_1 = {io_data_out_hi_hi_hi,io_data_out_hi_hi_hi,io_data_out_hi_hi_hi,io_data_out_hi_hi_hi,
    io_data_out_hi_hi_hi,io_data_out_hi_hi_hi,io_data_out_hi_hi_hi,io_data_out_hi_hi_hi}; // @[Cat.scala 30:58]
  wire [7:0] _io_data_out_T_2 = 8'h1b & _io_data_out_T_1; // @[GFMult.scala 13:42]
  wire [7:0] _io_data_out_T_3 = m[7:0] ^ _io_data_out_T_2; // @[GFMult.scala 13:24]
  wire  io_data_out_hi_hi_hi_1 = m[9]; // @[GFMult.scala 13:118]
  wire [7:0] _io_data_out_T_4 = {io_data_out_hi_hi_hi_1,io_data_out_hi_hi_hi_1,io_data_out_hi_hi_hi_1,
    io_data_out_hi_hi_hi_1,io_data_out_hi_hi_hi_1,io_data_out_hi_hi_hi_1,io_data_out_hi_hi_hi_1,io_data_out_hi_hi_hi_1}; // @[Cat.scala 30:58]
  wire [7:0] _io_data_out_T_5 = 8'h36 & _io_data_out_T_4; // @[GFMult.scala 13:110]
  wire [7:0] _io_data_out_T_6 = _io_data_out_T_3 ^ _io_data_out_T_5; // @[GFMult.scala 13:92]
  wire  io_data_out_hi_hi_hi_2 = m[10]; // @[GFMult.scala 13:187]
  wire [7:0] _io_data_out_T_7 = {io_data_out_hi_hi_hi_2,io_data_out_hi_hi_hi_2,io_data_out_hi_hi_hi_2,
    io_data_out_hi_hi_hi_2,io_data_out_hi_hi_hi_2,io_data_out_hi_hi_hi_2,io_data_out_hi_hi_hi_2,io_data_out_hi_hi_hi_2}; // @[Cat.scala 30:58]
  wire [7:0] _io_data_out_T_8 = 8'h6c & _io_data_out_T_7; // @[GFMult.scala 13:179]
  assign io_data_out = _io_data_out_T_6 ^ _io_data_out_T_8; // @[GFMult.scala 13:160]
endmodule
*/
module BS_MC(
  input  [127:0] io_data_in,
  output [127:0] io_data_out
);
  wire [127:0] bs_data_out_m_io_data_in; // @[BS_MC.scala 88:19]
  wire [127:0] bs_data_out_m_io_data_out; // @[BS_MC.scala 88:19]
  wire [7:0] k0_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k0_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k0_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k0_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k0_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k0_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k0_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k0_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k0_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k0_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k0_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k0_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k1_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k2_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k3_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k4_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k5_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k6_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k7_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k8_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k9_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k10_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k11_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k12_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k13_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k14_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_1_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_1_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_1_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_2_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_2_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_2_io_data_out; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_3_io_data_in_1; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_3_io_data_in_2; // @[GFMult.scala 18:19]
  wire [7:0] k15_a_3_io_data_out; // @[GFMult.scala 18:19]
  wire [127:0] bs_data_out = bs_data_out_m_io_data_out; // @[BS_MC.scala 45:25 BS_MC.scala 46:15]
  wire [7:0] _k0_T_2 = k0_a_io_data_out ^ k0_a_1_io_data_out; // @[BS_MC.scala 48:45]
  wire [7:0] _k0_T_4 = _k0_T_2 ^ k0_a_2_io_data_out; // @[BS_MC.scala 48:82]
  wire [7:0] k0 = _k0_T_4 ^ k0_a_3_io_data_out; // @[BS_MC.scala 48:120]
  wire [7:0] _k1_T_2 = k1_a_io_data_out ^ k1_a_1_io_data_out; // @[BS_MC.scala 49:45]
  wire [7:0] _k1_T_4 = _k1_T_2 ^ k1_a_2_io_data_out; // @[BS_MC.scala 49:82]
  wire [7:0] k1 = _k1_T_4 ^ k1_a_3_io_data_out; // @[BS_MC.scala 49:120]
  wire [7:0] _k2_T_2 = k2_a_io_data_out ^ k2_a_1_io_data_out; // @[BS_MC.scala 50:45]
  wire [7:0] _k2_T_4 = _k2_T_2 ^ k2_a_2_io_data_out; // @[BS_MC.scala 50:82]
  wire [7:0] k2 = _k2_T_4 ^ k2_a_3_io_data_out; // @[BS_MC.scala 50:120]
  wire [7:0] _k3_T_2 = k3_a_io_data_out ^ k3_a_1_io_data_out; // @[BS_MC.scala 51:45]
  wire [7:0] _k3_T_4 = _k3_T_2 ^ k3_a_2_io_data_out; // @[BS_MC.scala 51:82]
  wire [7:0] k3 = _k3_T_4 ^ k3_a_3_io_data_out; // @[BS_MC.scala 51:120]
  wire [7:0] _k4_T_2 = k4_a_io_data_out ^ k4_a_1_io_data_out; // @[BS_MC.scala 53:47]
  wire [7:0] _k4_T_4 = _k4_T_2 ^ k4_a_2_io_data_out; // @[BS_MC.scala 53:85]
  wire [7:0] k4 = _k4_T_4 ^ k4_a_3_io_data_out; // @[BS_MC.scala 53:123]
  wire [7:0] _k5_T_2 = k5_a_io_data_out ^ k5_a_1_io_data_out; // @[BS_MC.scala 54:47]
  wire [7:0] _k5_T_4 = _k5_T_2 ^ k5_a_2_io_data_out; // @[BS_MC.scala 54:85]
  wire [7:0] k5 = _k5_T_4 ^ k5_a_3_io_data_out; // @[BS_MC.scala 54:123]
  wire [7:0] _k6_T_2 = k6_a_io_data_out ^ k6_a_1_io_data_out; // @[BS_MC.scala 55:47]
  wire [7:0] _k6_T_4 = _k6_T_2 ^ k6_a_2_io_data_out; // @[BS_MC.scala 55:85]
  wire [7:0] k6 = _k6_T_4 ^ k6_a_3_io_data_out; // @[BS_MC.scala 55:123]
  wire [7:0] _k7_T_2 = k7_a_io_data_out ^ k7_a_1_io_data_out; // @[BS_MC.scala 56:47]
  wire [7:0] _k7_T_4 = _k7_T_2 ^ k7_a_2_io_data_out; // @[BS_MC.scala 56:85]
  wire [7:0] k7 = _k7_T_4 ^ k7_a_3_io_data_out; // @[BS_MC.scala 56:123]
  wire [7:0] _k8_T_2 = k8_a_io_data_out ^ k8_a_1_io_data_out; // @[BS_MC.scala 58:48]
  wire [7:0] _k8_T_4 = _k8_T_2 ^ k8_a_2_io_data_out; // @[BS_MC.scala 58:86]
  wire [7:0] k8 = _k8_T_4 ^ k8_a_3_io_data_out; // @[BS_MC.scala 58:124]
  wire [7:0] _k9_T_2 = k9_a_io_data_out ^ k9_a_1_io_data_out; // @[BS_MC.scala 59:48]
  wire [7:0] _k9_T_4 = _k9_T_2 ^ k9_a_2_io_data_out; // @[BS_MC.scala 59:86]
  wire [7:0] k9 = _k9_T_4 ^ k9_a_3_io_data_out; // @[BS_MC.scala 59:124]
  wire [7:0] _k10_T_2 = k10_a_io_data_out ^ k10_a_1_io_data_out; // @[BS_MC.scala 60:48]
  wire [7:0] _k10_T_4 = _k10_T_2 ^ k10_a_2_io_data_out; // @[BS_MC.scala 60:86]
  wire [7:0] k10 = _k10_T_4 ^ k10_a_3_io_data_out; // @[BS_MC.scala 60:124]
  wire [7:0] _k11_T_2 = k11_a_io_data_out ^ k11_a_1_io_data_out; // @[BS_MC.scala 61:48]
  wire [7:0] _k11_T_4 = _k11_T_2 ^ k11_a_2_io_data_out; // @[BS_MC.scala 61:86]
  wire [7:0] k11 = _k11_T_4 ^ k11_a_3_io_data_out; // @[BS_MC.scala 61:124]
  wire [7:0] _k12_T_2 = k12_a_io_data_out ^ k12_a_1_io_data_out; // @[BS_MC.scala 63:49]
  wire [7:0] _k12_T_4 = _k12_T_2 ^ k12_a_2_io_data_out; // @[BS_MC.scala 63:89]
  wire [7:0] k12 = _k12_T_4 ^ k12_a_3_io_data_out; // @[BS_MC.scala 63:129]
  wire [7:0] _k13_T_2 = k13_a_io_data_out ^ k13_a_1_io_data_out; // @[BS_MC.scala 64:49]
  wire [7:0] _k13_T_4 = _k13_T_2 ^ k13_a_2_io_data_out; // @[BS_MC.scala 64:89]
  wire [7:0] k13 = _k13_T_4 ^ k13_a_3_io_data_out; // @[BS_MC.scala 64:129]
  wire [7:0] _k14_T_2 = k14_a_io_data_out ^ k14_a_1_io_data_out; // @[BS_MC.scala 65:49]
  wire [7:0] _k14_T_4 = _k14_T_2 ^ k14_a_2_io_data_out; // @[BS_MC.scala 65:89]
  wire [7:0] k14 = _k14_T_4 ^ k14_a_3_io_data_out; // @[BS_MC.scala 65:129]
  wire [7:0] _k15_T_2 = k15_a_io_data_out ^ k15_a_1_io_data_out; // @[BS_MC.scala 66:49]
  wire [7:0] _k15_T_4 = _k15_T_2 ^ k15_a_2_io_data_out; // @[BS_MC.scala 66:89]
  wire [7:0] k15 = _k15_T_4 ^ k15_a_3_io_data_out; // @[BS_MC.scala 66:129]
  wire [63:0] io_data_out_lo = {k7,k6,k5,k4,k3,k2,k1,k0}; // @[Cat.scala 30:58]
  wire [63:0] io_data_out_hi = {k15,k14,k13,k12,k11,k10,k9,k8}; // @[Cat.scala 30:58]
  BS bs_data_out_m ( // @[BS_MC.scala 88:19]
    .io_data_in(bs_data_out_m_io_data_in),
    .io_data_out(bs_data_out_m_io_data_out)
  );
  GFMult k0_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k0_a_io_data_in_1),
    .io_data_in_2(k0_a_io_data_in_2),
    .io_data_out(k0_a_io_data_out)
  );
  GFMult k0_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k0_a_1_io_data_in_1),
    .io_data_in_2(k0_a_1_io_data_in_2),
    .io_data_out(k0_a_1_io_data_out)
  );
  GFMult k0_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k0_a_2_io_data_in_1),
    .io_data_in_2(k0_a_2_io_data_in_2),
    .io_data_out(k0_a_2_io_data_out)
  );
  GFMult k0_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k0_a_3_io_data_in_1),
    .io_data_in_2(k0_a_3_io_data_in_2),
    .io_data_out(k0_a_3_io_data_out)
  );
  GFMult k1_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k1_a_io_data_in_1),
    .io_data_in_2(k1_a_io_data_in_2),
    .io_data_out(k1_a_io_data_out)
  );
  GFMult k1_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k1_a_1_io_data_in_1),
    .io_data_in_2(k1_a_1_io_data_in_2),
    .io_data_out(k1_a_1_io_data_out)
  );
  GFMult k1_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k1_a_2_io_data_in_1),
    .io_data_in_2(k1_a_2_io_data_in_2),
    .io_data_out(k1_a_2_io_data_out)
  );
  GFMult k1_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k1_a_3_io_data_in_1),
    .io_data_in_2(k1_a_3_io_data_in_2),
    .io_data_out(k1_a_3_io_data_out)
  );
  GFMult k2_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k2_a_io_data_in_1),
    .io_data_in_2(k2_a_io_data_in_2),
    .io_data_out(k2_a_io_data_out)
  );
  GFMult k2_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k2_a_1_io_data_in_1),
    .io_data_in_2(k2_a_1_io_data_in_2),
    .io_data_out(k2_a_1_io_data_out)
  );
  GFMult k2_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k2_a_2_io_data_in_1),
    .io_data_in_2(k2_a_2_io_data_in_2),
    .io_data_out(k2_a_2_io_data_out)
  );
  GFMult k2_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k2_a_3_io_data_in_1),
    .io_data_in_2(k2_a_3_io_data_in_2),
    .io_data_out(k2_a_3_io_data_out)
  );
  GFMult k3_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k3_a_io_data_in_1),
    .io_data_in_2(k3_a_io_data_in_2),
    .io_data_out(k3_a_io_data_out)
  );
  GFMult k3_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k3_a_1_io_data_in_1),
    .io_data_in_2(k3_a_1_io_data_in_2),
    .io_data_out(k3_a_1_io_data_out)
  );
  GFMult k3_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k3_a_2_io_data_in_1),
    .io_data_in_2(k3_a_2_io_data_in_2),
    .io_data_out(k3_a_2_io_data_out)
  );
  GFMult k3_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k3_a_3_io_data_in_1),
    .io_data_in_2(k3_a_3_io_data_in_2),
    .io_data_out(k3_a_3_io_data_out)
  );
  GFMult k4_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k4_a_io_data_in_1),
    .io_data_in_2(k4_a_io_data_in_2),
    .io_data_out(k4_a_io_data_out)
  );
  GFMult k4_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k4_a_1_io_data_in_1),
    .io_data_in_2(k4_a_1_io_data_in_2),
    .io_data_out(k4_a_1_io_data_out)
  );
  GFMult k4_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k4_a_2_io_data_in_1),
    .io_data_in_2(k4_a_2_io_data_in_2),
    .io_data_out(k4_a_2_io_data_out)
  );
  GFMult k4_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k4_a_3_io_data_in_1),
    .io_data_in_2(k4_a_3_io_data_in_2),
    .io_data_out(k4_a_3_io_data_out)
  );
  GFMult k5_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k5_a_io_data_in_1),
    .io_data_in_2(k5_a_io_data_in_2),
    .io_data_out(k5_a_io_data_out)
  );
  GFMult k5_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k5_a_1_io_data_in_1),
    .io_data_in_2(k5_a_1_io_data_in_2),
    .io_data_out(k5_a_1_io_data_out)
  );
  GFMult k5_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k5_a_2_io_data_in_1),
    .io_data_in_2(k5_a_2_io_data_in_2),
    .io_data_out(k5_a_2_io_data_out)
  );
  GFMult k5_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k5_a_3_io_data_in_1),
    .io_data_in_2(k5_a_3_io_data_in_2),
    .io_data_out(k5_a_3_io_data_out)
  );
  GFMult k6_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k6_a_io_data_in_1),
    .io_data_in_2(k6_a_io_data_in_2),
    .io_data_out(k6_a_io_data_out)
  );
  GFMult k6_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k6_a_1_io_data_in_1),
    .io_data_in_2(k6_a_1_io_data_in_2),
    .io_data_out(k6_a_1_io_data_out)
  );
  GFMult k6_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k6_a_2_io_data_in_1),
    .io_data_in_2(k6_a_2_io_data_in_2),
    .io_data_out(k6_a_2_io_data_out)
  );
  GFMult k6_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k6_a_3_io_data_in_1),
    .io_data_in_2(k6_a_3_io_data_in_2),
    .io_data_out(k6_a_3_io_data_out)
  );
  GFMult k7_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k7_a_io_data_in_1),
    .io_data_in_2(k7_a_io_data_in_2),
    .io_data_out(k7_a_io_data_out)
  );
  GFMult k7_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k7_a_1_io_data_in_1),
    .io_data_in_2(k7_a_1_io_data_in_2),
    .io_data_out(k7_a_1_io_data_out)
  );
  GFMult k7_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k7_a_2_io_data_in_1),
    .io_data_in_2(k7_a_2_io_data_in_2),
    .io_data_out(k7_a_2_io_data_out)
  );
  GFMult k7_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k7_a_3_io_data_in_1),
    .io_data_in_2(k7_a_3_io_data_in_2),
    .io_data_out(k7_a_3_io_data_out)
  );
  GFMult k8_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k8_a_io_data_in_1),
    .io_data_in_2(k8_a_io_data_in_2),
    .io_data_out(k8_a_io_data_out)
  );
  GFMult k8_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k8_a_1_io_data_in_1),
    .io_data_in_2(k8_a_1_io_data_in_2),
    .io_data_out(k8_a_1_io_data_out)
  );
  GFMult k8_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k8_a_2_io_data_in_1),
    .io_data_in_2(k8_a_2_io_data_in_2),
    .io_data_out(k8_a_2_io_data_out)
  );
  GFMult k8_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k8_a_3_io_data_in_1),
    .io_data_in_2(k8_a_3_io_data_in_2),
    .io_data_out(k8_a_3_io_data_out)
  );
  GFMult k9_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k9_a_io_data_in_1),
    .io_data_in_2(k9_a_io_data_in_2),
    .io_data_out(k9_a_io_data_out)
  );
  GFMult k9_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k9_a_1_io_data_in_1),
    .io_data_in_2(k9_a_1_io_data_in_2),
    .io_data_out(k9_a_1_io_data_out)
  );
  GFMult k9_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k9_a_2_io_data_in_1),
    .io_data_in_2(k9_a_2_io_data_in_2),
    .io_data_out(k9_a_2_io_data_out)
  );
  GFMult k9_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k9_a_3_io_data_in_1),
    .io_data_in_2(k9_a_3_io_data_in_2),
    .io_data_out(k9_a_3_io_data_out)
  );
  GFMult k10_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k10_a_io_data_in_1),
    .io_data_in_2(k10_a_io_data_in_2),
    .io_data_out(k10_a_io_data_out)
  );
  GFMult k10_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k10_a_1_io_data_in_1),
    .io_data_in_2(k10_a_1_io_data_in_2),
    .io_data_out(k10_a_1_io_data_out)
  );
  GFMult k10_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k10_a_2_io_data_in_1),
    .io_data_in_2(k10_a_2_io_data_in_2),
    .io_data_out(k10_a_2_io_data_out)
  );
  GFMult k10_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k10_a_3_io_data_in_1),
    .io_data_in_2(k10_a_3_io_data_in_2),
    .io_data_out(k10_a_3_io_data_out)
  );
  GFMult k11_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k11_a_io_data_in_1),
    .io_data_in_2(k11_a_io_data_in_2),
    .io_data_out(k11_a_io_data_out)
  );
  GFMult k11_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k11_a_1_io_data_in_1),
    .io_data_in_2(k11_a_1_io_data_in_2),
    .io_data_out(k11_a_1_io_data_out)
  );
  GFMult k11_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k11_a_2_io_data_in_1),
    .io_data_in_2(k11_a_2_io_data_in_2),
    .io_data_out(k11_a_2_io_data_out)
  );
  GFMult k11_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k11_a_3_io_data_in_1),
    .io_data_in_2(k11_a_3_io_data_in_2),
    .io_data_out(k11_a_3_io_data_out)
  );
  GFMult k12_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k12_a_io_data_in_1),
    .io_data_in_2(k12_a_io_data_in_2),
    .io_data_out(k12_a_io_data_out)
  );
  GFMult k12_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k12_a_1_io_data_in_1),
    .io_data_in_2(k12_a_1_io_data_in_2),
    .io_data_out(k12_a_1_io_data_out)
  );
  GFMult k12_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k12_a_2_io_data_in_1),
    .io_data_in_2(k12_a_2_io_data_in_2),
    .io_data_out(k12_a_2_io_data_out)
  );
  GFMult k12_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k12_a_3_io_data_in_1),
    .io_data_in_2(k12_a_3_io_data_in_2),
    .io_data_out(k12_a_3_io_data_out)
  );
  GFMult k13_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k13_a_io_data_in_1),
    .io_data_in_2(k13_a_io_data_in_2),
    .io_data_out(k13_a_io_data_out)
  );
  GFMult k13_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k13_a_1_io_data_in_1),
    .io_data_in_2(k13_a_1_io_data_in_2),
    .io_data_out(k13_a_1_io_data_out)
  );
  GFMult k13_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k13_a_2_io_data_in_1),
    .io_data_in_2(k13_a_2_io_data_in_2),
    .io_data_out(k13_a_2_io_data_out)
  );
  GFMult k13_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k13_a_3_io_data_in_1),
    .io_data_in_2(k13_a_3_io_data_in_2),
    .io_data_out(k13_a_3_io_data_out)
  );
  GFMult k14_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k14_a_io_data_in_1),
    .io_data_in_2(k14_a_io_data_in_2),
    .io_data_out(k14_a_io_data_out)
  );
  GFMult k14_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k14_a_1_io_data_in_1),
    .io_data_in_2(k14_a_1_io_data_in_2),
    .io_data_out(k14_a_1_io_data_out)
  );
  GFMult k14_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k14_a_2_io_data_in_1),
    .io_data_in_2(k14_a_2_io_data_in_2),
    .io_data_out(k14_a_2_io_data_out)
  );
  GFMult k14_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k14_a_3_io_data_in_1),
    .io_data_in_2(k14_a_3_io_data_in_2),
    .io_data_out(k14_a_3_io_data_out)
  );
  GFMult k15_a ( // @[GFMult.scala 18:19]
    .io_data_in_1(k15_a_io_data_in_1),
    .io_data_in_2(k15_a_io_data_in_2),
    .io_data_out(k15_a_io_data_out)
  );
  GFMult k15_a_1 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k15_a_1_io_data_in_1),
    .io_data_in_2(k15_a_1_io_data_in_2),
    .io_data_out(k15_a_1_io_data_out)
  );
  GFMult k15_a_2 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k15_a_2_io_data_in_1),
    .io_data_in_2(k15_a_2_io_data_in_2),
    .io_data_out(k15_a_2_io_data_out)
  );
  GFMult k15_a_3 ( // @[GFMult.scala 18:19]
    .io_data_in_1(k15_a_3_io_data_in_1),
    .io_data_in_2(k15_a_3_io_data_in_2),
    .io_data_out(k15_a_3_io_data_out)
  );
  assign io_data_out = {io_data_out_hi,io_data_out_lo}; // @[Cat.scala 30:58]
  assign bs_data_out_m_io_data_in = io_data_in; // @[BS_MC.scala 89:18]
  assign k0_a_io_data_in_1 = bs_data_out[7:0]; // @[BS_MC.scala 48:38]
  assign k0_a_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k0_a_1_io_data_in_1 = bs_data_out[15:8]; // @[BS_MC.scala 48:74]
  assign k0_a_1_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k0_a_2_io_data_in_1 = bs_data_out[23:16]; // @[BS_MC.scala 48:111]
  assign k0_a_2_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k0_a_3_io_data_in_1 = bs_data_out[31:24]; // @[BS_MC.scala 48:149]
  assign k0_a_3_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k1_a_io_data_in_1 = bs_data_out[7:0]; // @[BS_MC.scala 49:38]
  assign k1_a_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k1_a_1_io_data_in_1 = bs_data_out[15:8]; // @[BS_MC.scala 49:74]
  assign k1_a_1_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k1_a_2_io_data_in_1 = bs_data_out[23:16]; // @[BS_MC.scala 49:111]
  assign k1_a_2_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k1_a_3_io_data_in_1 = bs_data_out[31:24]; // @[BS_MC.scala 49:149]
  assign k1_a_3_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k2_a_io_data_in_1 = bs_data_out[7:0]; // @[BS_MC.scala 50:38]
  assign k2_a_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k2_a_1_io_data_in_1 = bs_data_out[15:8]; // @[BS_MC.scala 50:74]
  assign k2_a_1_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k2_a_2_io_data_in_1 = bs_data_out[23:16]; // @[BS_MC.scala 50:111]
  assign k2_a_2_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k2_a_3_io_data_in_1 = bs_data_out[31:24]; // @[BS_MC.scala 50:149]
  assign k2_a_3_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k3_a_io_data_in_1 = bs_data_out[7:0]; // @[BS_MC.scala 51:38]
  assign k3_a_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k3_a_1_io_data_in_1 = bs_data_out[15:8]; // @[BS_MC.scala 51:74]
  assign k3_a_1_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k3_a_2_io_data_in_1 = bs_data_out[23:16]; // @[BS_MC.scala 51:111]
  assign k3_a_2_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k3_a_3_io_data_in_1 = bs_data_out[31:24]; // @[BS_MC.scala 51:149]
  assign k3_a_3_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k4_a_io_data_in_1 = bs_data_out[39:32]; // @[BS_MC.scala 53:38]
  assign k4_a_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k4_a_1_io_data_in_1 = bs_data_out[47:40]; // @[BS_MC.scala 53:76]
  assign k4_a_1_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k4_a_2_io_data_in_1 = bs_data_out[55:48]; // @[BS_MC.scala 53:114]
  assign k4_a_2_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k4_a_3_io_data_in_1 = bs_data_out[63:56]; // @[BS_MC.scala 53:152]
  assign k4_a_3_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k5_a_io_data_in_1 = bs_data_out[39:32]; // @[BS_MC.scala 54:38]
  assign k5_a_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k5_a_1_io_data_in_1 = bs_data_out[47:40]; // @[BS_MC.scala 54:76]
  assign k5_a_1_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k5_a_2_io_data_in_1 = bs_data_out[55:48]; // @[BS_MC.scala 54:114]
  assign k5_a_2_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k5_a_3_io_data_in_1 = bs_data_out[63:56]; // @[BS_MC.scala 54:152]
  assign k5_a_3_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k6_a_io_data_in_1 = bs_data_out[39:32]; // @[BS_MC.scala 55:38]
  assign k6_a_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k6_a_1_io_data_in_1 = bs_data_out[47:40]; // @[BS_MC.scala 55:76]
  assign k6_a_1_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k6_a_2_io_data_in_1 = bs_data_out[55:48]; // @[BS_MC.scala 55:114]
  assign k6_a_2_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k6_a_3_io_data_in_1 = bs_data_out[63:56]; // @[BS_MC.scala 55:152]
  assign k6_a_3_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k7_a_io_data_in_1 = bs_data_out[39:32]; // @[BS_MC.scala 56:38]
  assign k7_a_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k7_a_1_io_data_in_1 = bs_data_out[47:40]; // @[BS_MC.scala 56:76]
  assign k7_a_1_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k7_a_2_io_data_in_1 = bs_data_out[55:48]; // @[BS_MC.scala 56:114]
  assign k7_a_2_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k7_a_3_io_data_in_1 = bs_data_out[63:56]; // @[BS_MC.scala 56:152]
  assign k7_a_3_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k8_a_io_data_in_1 = bs_data_out[71:64]; // @[BS_MC.scala 58:39]
  assign k8_a_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k8_a_1_io_data_in_1 = bs_data_out[79:72]; // @[BS_MC.scala 58:77]
  assign k8_a_1_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k8_a_2_io_data_in_1 = bs_data_out[87:80]; // @[BS_MC.scala 58:115]
  assign k8_a_2_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k8_a_3_io_data_in_1 = bs_data_out[95:88]; // @[BS_MC.scala 58:153]
  assign k8_a_3_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k9_a_io_data_in_1 = bs_data_out[71:64]; // @[BS_MC.scala 59:39]
  assign k9_a_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k9_a_1_io_data_in_1 = bs_data_out[79:72]; // @[BS_MC.scala 59:77]
  assign k9_a_1_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k9_a_2_io_data_in_1 = bs_data_out[87:80]; // @[BS_MC.scala 59:115]
  assign k9_a_2_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k9_a_3_io_data_in_1 = bs_data_out[95:88]; // @[BS_MC.scala 59:153]
  assign k9_a_3_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k10_a_io_data_in_1 = bs_data_out[71:64]; // @[BS_MC.scala 60:39]
  assign k10_a_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k10_a_1_io_data_in_1 = bs_data_out[79:72]; // @[BS_MC.scala 60:77]
  assign k10_a_1_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k10_a_2_io_data_in_1 = bs_data_out[87:80]; // @[BS_MC.scala 60:115]
  assign k10_a_2_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k10_a_3_io_data_in_1 = bs_data_out[95:88]; // @[BS_MC.scala 60:153]
  assign k10_a_3_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k11_a_io_data_in_1 = bs_data_out[71:64]; // @[BS_MC.scala 61:39]
  assign k11_a_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k11_a_1_io_data_in_1 = bs_data_out[79:72]; // @[BS_MC.scala 61:77]
  assign k11_a_1_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k11_a_2_io_data_in_1 = bs_data_out[87:80]; // @[BS_MC.scala 61:115]
  assign k11_a_2_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k11_a_3_io_data_in_1 = bs_data_out[95:88]; // @[BS_MC.scala 61:153]
  assign k11_a_3_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k12_a_io_data_in_1 = bs_data_out[103:96]; // @[BS_MC.scala 63:39]
  assign k12_a_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k12_a_1_io_data_in_1 = bs_data_out[111:104]; // @[BS_MC.scala 63:78]
  assign k12_a_1_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k12_a_2_io_data_in_1 = bs_data_out[119:112]; // @[BS_MC.scala 63:118]
  assign k12_a_2_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k12_a_3_io_data_in_1 = bs_data_out[127:120]; // @[BS_MC.scala 63:158]
  assign k12_a_3_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k13_a_io_data_in_1 = bs_data_out[103:96]; // @[BS_MC.scala 64:39]
  assign k13_a_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k13_a_1_io_data_in_1 = bs_data_out[111:104]; // @[BS_MC.scala 64:78]
  assign k13_a_1_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k13_a_2_io_data_in_1 = bs_data_out[119:112]; // @[BS_MC.scala 64:118]
  assign k13_a_2_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k13_a_3_io_data_in_1 = bs_data_out[127:120]; // @[BS_MC.scala 64:158]
  assign k13_a_3_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k14_a_io_data_in_1 = bs_data_out[103:96]; // @[BS_MC.scala 65:39]
  assign k14_a_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k14_a_1_io_data_in_1 = bs_data_out[111:104]; // @[BS_MC.scala 65:78]
  assign k14_a_1_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k14_a_2_io_data_in_1 = bs_data_out[119:112]; // @[BS_MC.scala 65:118]
  assign k14_a_2_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
  assign k14_a_3_io_data_in_1 = bs_data_out[127:120]; // @[BS_MC.scala 65:158]
  assign k14_a_3_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k15_a_io_data_in_1 = bs_data_out[103:96]; // @[BS_MC.scala 66:39]
  assign k15_a_io_data_in_2 = 8'h3; // @[GFMult.scala 20:20]
  assign k15_a_1_io_data_in_1 = bs_data_out[111:104]; // @[BS_MC.scala 66:78]
  assign k15_a_1_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k15_a_2_io_data_in_1 = bs_data_out[119:112]; // @[BS_MC.scala 66:118]
  assign k15_a_2_io_data_in_2 = 8'h1; // @[GFMult.scala 20:20]
  assign k15_a_3_io_data_in_1 = bs_data_out[127:120]; // @[BS_MC.scala 66:158]
  assign k15_a_3_io_data_in_2 = 8'h2; // @[GFMult.scala 20:20]
endmodule
module AES128(
  input          clock,
  input          reset,
  input  [127:0] io_data_in,
  input  [127:0] io_key_in,
  output [127:0] io_data_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] round0_data_out_a_io_data_in_1; // @[XOR32.scala 22:19]
  wire [127:0] round0_data_out_a_io_data_in_2; // @[XOR32.scala 22:19]
  wire [127:0] round0_data_out_a_io_data_out; // @[XOR32.scala 22:19]
  wire [31:0] w4_g_io_data_in; // @[G_func.scala 14:19]
  wire [7:0] w4_g_io_rc_in; // @[G_func.scala 14:19]
  wire [31:0] w4_g_io_data_out; // @[G_func.scala 14:19]
  wire [31:0] w4_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w4_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w4_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w5_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w5_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w5_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w6_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w6_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w6_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w7_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w7_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w7_a_io_data_out; // @[XOR32.scala 9:19]
  wire [127:0] data_c1_SR_io_data_in; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c1_SR_io_data_out; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c1_m_io_data_in; // @[BS_MC.scala 72:19]
  wire [127:0] data_c1_m_io_data_out; // @[BS_MC.scala 72:19]
  wire [127:0] round1_data_out_a_io_data_in_1; // @[XOR32.scala 22:19]
  wire [127:0] round1_data_out_a_io_data_in_2; // @[XOR32.scala 22:19]
  wire [127:0] round1_data_out_a_io_data_out; // @[XOR32.scala 22:19]
  wire [31:0] w8_g_io_data_in; // @[G_func.scala 14:19]
  wire [7:0] w8_g_io_rc_in; // @[G_func.scala 14:19]
  wire [31:0] w8_g_io_data_out; // @[G_func.scala 14:19]
  wire [31:0] w8_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w8_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w8_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w9_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w9_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w9_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w10_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w10_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w10_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w11_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w11_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w11_a_io_data_out; // @[XOR32.scala 9:19]
  wire [127:0] data_c2_SR_io_data_in; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c2_SR_io_data_out; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c2_m_io_data_in; // @[BS_MC.scala 72:19]
  wire [127:0] data_c2_m_io_data_out; // @[BS_MC.scala 72:19]
  wire [127:0] round2_data_out_a_io_data_in_1; // @[XOR32.scala 22:19]
  wire [127:0] round2_data_out_a_io_data_in_2; // @[XOR32.scala 22:19]
  wire [127:0] round2_data_out_a_io_data_out; // @[XOR32.scala 22:19]
  wire [31:0] w12_g_io_data_in; // @[G_func.scala 14:19]
  wire [7:0] w12_g_io_rc_in; // @[G_func.scala 14:19]
  wire [31:0] w12_g_io_data_out; // @[G_func.scala 14:19]
  wire [31:0] w12_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w12_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w12_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w13_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w13_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w13_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w14_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w14_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w14_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w15_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w15_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w15_a_io_data_out; // @[XOR32.scala 9:19]
  wire [127:0] data_c3_SR_io_data_in; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c3_SR_io_data_out; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c3_m_io_data_in; // @[BS_MC.scala 72:19]
  wire [127:0] data_c3_m_io_data_out; // @[BS_MC.scala 72:19]
  wire [127:0] round3_data_out_a_io_data_in_1; // @[XOR32.scala 22:19]
  wire [127:0] round3_data_out_a_io_data_in_2; // @[XOR32.scala 22:19]
  wire [127:0] round3_data_out_a_io_data_out; // @[XOR32.scala 22:19]
  wire [31:0] w16_g_io_data_in; // @[G_func.scala 14:19]
  wire [7:0] w16_g_io_rc_in; // @[G_func.scala 14:19]
  wire [31:0] w16_g_io_data_out; // @[G_func.scala 14:19]
  wire [31:0] w16_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w16_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w16_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w17_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w17_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w17_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w18_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w18_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w18_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w19_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w19_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w19_a_io_data_out; // @[XOR32.scala 9:19]
  wire [127:0] data_c4_SR_io_data_in; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c4_SR_io_data_out; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c4_m_io_data_in; // @[BS_MC.scala 72:19]
  wire [127:0] data_c4_m_io_data_out; // @[BS_MC.scala 72:19]
  wire [127:0] round4_data_out_a_io_data_in_1; // @[XOR32.scala 22:19]
  wire [127:0] round4_data_out_a_io_data_in_2; // @[XOR32.scala 22:19]
  wire [127:0] round4_data_out_a_io_data_out; // @[XOR32.scala 22:19]
  wire [31:0] w20_g_io_data_in; // @[G_func.scala 14:19]
  wire [7:0] w20_g_io_rc_in; // @[G_func.scala 14:19]
  wire [31:0] w20_g_io_data_out; // @[G_func.scala 14:19]
  wire [31:0] w20_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w20_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w20_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w21_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w21_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w21_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w22_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w22_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w22_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w23_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w23_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w23_a_io_data_out; // @[XOR32.scala 9:19]
  wire [127:0] data_c5_SR_io_data_in; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c5_SR_io_data_out; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c5_m_io_data_in; // @[BS_MC.scala 72:19]
  wire [127:0] data_c5_m_io_data_out; // @[BS_MC.scala 72:19]
  wire [127:0] round5_data_out_a_io_data_in_1; // @[XOR32.scala 22:19]
  wire [127:0] round5_data_out_a_io_data_in_2; // @[XOR32.scala 22:19]
  wire [127:0] round5_data_out_a_io_data_out; // @[XOR32.scala 22:19]
  wire [31:0] w24_g_io_data_in; // @[G_func.scala 14:19]
  wire [7:0] w24_g_io_rc_in; // @[G_func.scala 14:19]
  wire [31:0] w24_g_io_data_out; // @[G_func.scala 14:19]
  wire [31:0] w24_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w24_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w24_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w25_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w25_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w25_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w26_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w26_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w26_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w27_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w27_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w27_a_io_data_out; // @[XOR32.scala 9:19]
  wire [127:0] data_c6_SR_io_data_in; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c6_SR_io_data_out; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c6_m_io_data_in; // @[BS_MC.scala 72:19]
  wire [127:0] data_c6_m_io_data_out; // @[BS_MC.scala 72:19]
  wire [127:0] round6_data_out_a_io_data_in_1; // @[XOR32.scala 22:19]
  wire [127:0] round6_data_out_a_io_data_in_2; // @[XOR32.scala 22:19]
  wire [127:0] round6_data_out_a_io_data_out; // @[XOR32.scala 22:19]
  wire [31:0] w28_g_io_data_in; // @[G_func.scala 14:19]
  wire [7:0] w28_g_io_rc_in; // @[G_func.scala 14:19]
  wire [31:0] w28_g_io_data_out; // @[G_func.scala 14:19]
  wire [31:0] w28_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w28_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w28_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w29_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w29_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w29_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w30_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w30_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w30_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w31_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w31_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w31_a_io_data_out; // @[XOR32.scala 9:19]
  wire [127:0] data_c7_SR_io_data_in; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c7_SR_io_data_out; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c7_m_io_data_in; // @[BS_MC.scala 72:19]
  wire [127:0] data_c7_m_io_data_out; // @[BS_MC.scala 72:19]
  wire [127:0] round7_data_out_a_io_data_in_1; // @[XOR32.scala 22:19]
  wire [127:0] round7_data_out_a_io_data_in_2; // @[XOR32.scala 22:19]
  wire [127:0] round7_data_out_a_io_data_out; // @[XOR32.scala 22:19]
  wire [31:0] w32_g_io_data_in; // @[G_func.scala 14:19]
  wire [7:0] w32_g_io_rc_in; // @[G_func.scala 14:19]
  wire [31:0] w32_g_io_data_out; // @[G_func.scala 14:19]
  wire [31:0] w32_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w32_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w32_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w33_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w33_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w33_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w34_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w34_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w34_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w35_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w35_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w35_a_io_data_out; // @[XOR32.scala 9:19]
  wire [127:0] data_c8_SR_io_data_in; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c8_SR_io_data_out; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c8_m_io_data_in; // @[BS_MC.scala 72:19]
  wire [127:0] data_c8_m_io_data_out; // @[BS_MC.scala 72:19]
  wire [127:0] round8_data_out_a_io_data_in_1; // @[XOR32.scala 22:19]
  wire [127:0] round8_data_out_a_io_data_in_2; // @[XOR32.scala 22:19]
  wire [127:0] round8_data_out_a_io_data_out; // @[XOR32.scala 22:19]
  wire [31:0] w36_g_io_data_in; // @[G_func.scala 14:19]
  wire [7:0] w36_g_io_rc_in; // @[G_func.scala 14:19]
  wire [31:0] w36_g_io_data_out; // @[G_func.scala 14:19]
  wire [31:0] w36_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w36_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w36_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w37_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w37_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w37_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w38_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w38_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w38_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w39_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w39_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w39_a_io_data_out; // @[XOR32.scala 9:19]
  wire [127:0] data_c9_SR_io_data_in; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c9_SR_io_data_out; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c9_m_io_data_in; // @[BS_MC.scala 72:19]
  wire [127:0] data_c9_m_io_data_out; // @[BS_MC.scala 72:19]
  wire [127:0] round9_data_out_a_io_data_in_1; // @[XOR32.scala 22:19]
  wire [127:0] round9_data_out_a_io_data_in_2; // @[XOR32.scala 22:19]
  wire [127:0] round9_data_out_a_io_data_out; // @[XOR32.scala 22:19]
  wire [31:0] w40_g_io_data_in; // @[G_func.scala 14:19]
  wire [7:0] w40_g_io_rc_in; // @[G_func.scala 14:19]
  wire [31:0] w40_g_io_data_out; // @[G_func.scala 14:19]
  wire [31:0] w40_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w40_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w40_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w41_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w41_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w41_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w42_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w42_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w42_a_io_data_out; // @[XOR32.scala 9:19]
  wire [31:0] w43_a_io_data_in_1; // @[XOR32.scala 9:19]
  wire [31:0] w43_a_io_data_in_2; // @[XOR32.scala 9:19]
  wire [31:0] w43_a_io_data_out; // @[XOR32.scala 9:19]
  wire [127:0] data_c10_SR_io_data_in; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c10_SR_io_data_out; // @[ShiftRows.scala 14:20]
  wire [127:0] data_c10_m_io_data_in; // @[BS_MC.scala 88:19]
  wire [127:0] data_c10_m_io_data_out; // @[BS_MC.scala 88:19]
  wire [127:0] round10_data_out_a_io_data_in_1; // @[XOR32.scala 22:19]
  wire [127:0] round10_data_out_a_io_data_in_2; // @[XOR32.scala 22:19]
  wire [127:0] round10_data_out_a_io_data_out; // @[XOR32.scala 22:19]
  reg [127:0] data_r0; // @[AES128.scala 9:20]
  reg [127:0] key_r0; // @[AES128.scala 10:19]
  reg [127:0] data_r1; // @[AES128.scala 21:20]
  reg [127:0] key_r1; // @[AES128.scala 22:19]
  wire [31:0] w5 = w5_a_io_data_out; // @[AES128.scala 24:16 AES128.scala 30:6]
  wire [31:0] w4 = w4_a_io_data_out; // @[AES128.scala 23:16 AES128.scala 29:6]
  wire [31:0] w7 = w7_a_io_data_out; // @[AES128.scala 26:16 AES128.scala 32:6]
  wire [31:0] w6 = w6_a_io_data_out; // @[AES128.scala 25:16 AES128.scala 31:6]
  wire [127:0] _key_r1_T = {w7,w6,w5,w4}; // @[Cat.scala 30:58]
  wire [127:0] data_c1 = data_c1_m_io_data_out; // @[AES128.scala 27:21 AES128.scala 33:11]
  reg [127:0] data_r2; // @[AES128.scala 43:20]
  reg [127:0] key_r2; // @[AES128.scala 44:19]
  wire [31:0] w9 = w9_a_io_data_out; // @[AES128.scala 46:16 AES128.scala 52:6]
  wire [31:0] w8 = w8_a_io_data_out; // @[AES128.scala 45:16 AES128.scala 51:6]
  wire [31:0] w11 = w11_a_io_data_out; // @[AES128.scala 48:17 AES128.scala 54:7]
  wire [31:0] w10 = w10_a_io_data_out; // @[AES128.scala 47:17 AES128.scala 53:7]
  wire [127:0] _key_r2_T = {w11,w10,w9,w8}; // @[Cat.scala 30:58]
  wire [127:0] data_c2 = data_c2_m_io_data_out; // @[AES128.scala 49:21 AES128.scala 55:11]
  reg [127:0] data_r3; // @[AES128.scala 65:20]
  reg [127:0] key_r3; // @[AES128.scala 66:19]
  wire [31:0] w13 = w13_a_io_data_out; // @[AES128.scala 68:17 AES128.scala 74:7]
  wire [31:0] w12 = w12_a_io_data_out; // @[AES128.scala 67:17 AES128.scala 73:7]
  wire [31:0] w15 = w15_a_io_data_out; // @[AES128.scala 70:17 AES128.scala 76:7]
  wire [31:0] w14 = w14_a_io_data_out; // @[AES128.scala 69:17 AES128.scala 75:7]
  wire [127:0] _key_r3_T = {w15,w14,w13,w12}; // @[Cat.scala 30:58]
  wire [127:0] data_c3 = data_c3_m_io_data_out; // @[AES128.scala 71:21 AES128.scala 77:11]
  reg [127:0] data_r4; // @[AES128.scala 87:20]
  reg [127:0] key_r4; // @[AES128.scala 88:19]
  wire [31:0] w17 = w17_a_io_data_out; // @[AES128.scala 90:17 AES128.scala 96:7]
  wire [31:0] w16 = w16_a_io_data_out; // @[AES128.scala 89:17 AES128.scala 95:7]
  wire [31:0] w19 = w19_a_io_data_out; // @[AES128.scala 92:17 AES128.scala 98:7]
  wire [31:0] w18 = w18_a_io_data_out; // @[AES128.scala 91:17 AES128.scala 97:7]
  wire [127:0] _key_r4_T = {w19,w18,w17,w16}; // @[Cat.scala 30:58]
  wire [127:0] data_c4 = data_c4_m_io_data_out; // @[AES128.scala 93:21 AES128.scala 99:11]
  reg [127:0] data_r5; // @[AES128.scala 109:20]
  reg [127:0] key_r5; // @[AES128.scala 110:19]
  wire [31:0] w21 = w21_a_io_data_out; // @[AES128.scala 112:17 AES128.scala 118:7]
  wire [31:0] w20 = w20_a_io_data_out; // @[AES128.scala 111:17 AES128.scala 117:7]
  wire [31:0] w23 = w23_a_io_data_out; // @[AES128.scala 114:17 AES128.scala 120:7]
  wire [31:0] w22 = w22_a_io_data_out; // @[AES128.scala 113:17 AES128.scala 119:7]
  wire [127:0] _key_r5_T = {w23,w22,w21,w20}; // @[Cat.scala 30:58]
  wire [127:0] data_c5 = data_c5_m_io_data_out; // @[AES128.scala 115:21 AES128.scala 121:11]
  reg [127:0] data_r6; // @[AES128.scala 131:20]
  reg [127:0] key_r6; // @[AES128.scala 132:19]
  wire [31:0] w25 = w25_a_io_data_out; // @[AES128.scala 134:17 AES128.scala 140:7]
  wire [31:0] w24 = w24_a_io_data_out; // @[AES128.scala 133:17 AES128.scala 139:7]
  wire [31:0] w27 = w27_a_io_data_out; // @[AES128.scala 136:17 AES128.scala 142:7]
  wire [31:0] w26 = w26_a_io_data_out; // @[AES128.scala 135:17 AES128.scala 141:7]
  wire [127:0] _key_r6_T = {w27,w26,w25,w24}; // @[Cat.scala 30:58]
  wire [127:0] data_c6 = data_c6_m_io_data_out; // @[AES128.scala 137:21 AES128.scala 143:11]
  reg [127:0] data_r7; // @[AES128.scala 153:20]
  reg [127:0] key_r7; // @[AES128.scala 154:19]
  wire [31:0] w29 = w29_a_io_data_out; // @[AES128.scala 156:17 AES128.scala 162:7]
  wire [31:0] w28 = w28_a_io_data_out; // @[AES128.scala 155:17 AES128.scala 161:7]
  wire [31:0] w31 = w31_a_io_data_out; // @[AES128.scala 158:17 AES128.scala 164:7]
  wire [31:0] w30 = w30_a_io_data_out; // @[AES128.scala 157:17 AES128.scala 163:7]
  wire [127:0] _key_r7_T = {w31,w30,w29,w28}; // @[Cat.scala 30:58]
  wire [127:0] data_c7 = data_c7_m_io_data_out; // @[AES128.scala 159:21 AES128.scala 165:11]
  reg [127:0] data_r8; // @[AES128.scala 175:20]
  reg [127:0] key_r8; // @[AES128.scala 176:19]
  wire [31:0] w33 = w33_a_io_data_out; // @[AES128.scala 178:17 AES128.scala 184:7]
  wire [31:0] w32 = w32_a_io_data_out; // @[AES128.scala 177:17 AES128.scala 183:7]
  wire [31:0] w35 = w35_a_io_data_out; // @[AES128.scala 180:17 AES128.scala 186:7]
  wire [31:0] w34 = w34_a_io_data_out; // @[AES128.scala 179:17 AES128.scala 185:7]
  wire [127:0] _key_r8_T = {w35,w34,w33,w32}; // @[Cat.scala 30:58]
  wire [127:0] data_c8 = data_c8_m_io_data_out; // @[AES128.scala 181:21 AES128.scala 187:11]
  reg [127:0] data_r9; // @[AES128.scala 197:20]
  reg [127:0] key_r9; // @[AES128.scala 198:19]
  wire [31:0] w37 = w37_a_io_data_out; // @[AES128.scala 200:17 AES128.scala 206:7]
  wire [31:0] w36 = w36_a_io_data_out; // @[AES128.scala 199:17 AES128.scala 205:7]
  wire [31:0] w39 = w39_a_io_data_out; // @[AES128.scala 202:17 AES128.scala 208:7]
  wire [31:0] w38 = w38_a_io_data_out; // @[AES128.scala 201:17 AES128.scala 207:7]
  wire [127:0] _key_r9_T = {w39,w38,w37,w36}; // @[Cat.scala 30:58]
  wire [127:0] data_c9 = data_c9_m_io_data_out; // @[AES128.scala 203:21 AES128.scala 209:11]
  reg [127:0] data_r10; // @[AES128.scala 219:21]
  reg [127:0] key_r10; // @[AES128.scala 220:20]
  wire [31:0] w41 = w41_a_io_data_out; // @[AES128.scala 222:17 AES128.scala 228:7]
  wire [31:0] w40 = w40_a_io_data_out; // @[AES128.scala 221:17 AES128.scala 227:7]
  wire [31:0] w43 = w43_a_io_data_out; // @[AES128.scala 224:17 AES128.scala 230:7]
  wire [31:0] w42 = w42_a_io_data_out; // @[AES128.scala 223:17 AES128.scala 229:7]
  wire [127:0] _key_r10_T = {w43,w42,w41,w40}; // @[Cat.scala 30:58]
  wire [127:0] data_c10 = data_c10_m_io_data_out; // @[AES128.scala 225:22 AES128.scala 231:12]
  XOR128 round0_data_out_a ( // @[XOR32.scala 22:19]
    .io_data_in_1(round0_data_out_a_io_data_in_1),
    .io_data_in_2(round0_data_out_a_io_data_in_2),
    .io_data_out(round0_data_out_a_io_data_out)
  );
  G_func w4_g ( // @[G_func.scala 14:19]
    .io_data_in(w4_g_io_data_in),
    .io_rc_in(w4_g_io_rc_in),
    .io_data_out(w4_g_io_data_out)
  );
  XOR32 w4_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w4_a_io_data_in_1),
    .io_data_in_2(w4_a_io_data_in_2),
    .io_data_out(w4_a_io_data_out)
  );
  XOR32 w5_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w5_a_io_data_in_1),
    .io_data_in_2(w5_a_io_data_in_2),
    .io_data_out(w5_a_io_data_out)
  );
  XOR32 w6_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w6_a_io_data_in_1),
    .io_data_in_2(w6_a_io_data_in_2),
    .io_data_out(w6_a_io_data_out)
  );
  XOR32 w7_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w7_a_io_data_in_1),
    .io_data_in_2(w7_a_io_data_in_2),
    .io_data_out(w7_a_io_data_out)
  );
  ShiftRows data_c1_SR ( // @[ShiftRows.scala 14:20]
    .io_data_in(data_c1_SR_io_data_in),
    .io_data_out(data_c1_SR_io_data_out)
  );
  BS_MC data_c1_m ( // @[BS_MC.scala 72:19]
    .io_data_in(data_c1_m_io_data_in),
    .io_data_out(data_c1_m_io_data_out)
  );
  XOR128 round1_data_out_a ( // @[XOR32.scala 22:19]
    .io_data_in_1(round1_data_out_a_io_data_in_1),
    .io_data_in_2(round1_data_out_a_io_data_in_2),
    .io_data_out(round1_data_out_a_io_data_out)
  );
  G_func w8_g ( // @[G_func.scala 14:19]
    .io_data_in(w8_g_io_data_in),
    .io_rc_in(w8_g_io_rc_in),
    .io_data_out(w8_g_io_data_out)
  );
  XOR32 w8_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w8_a_io_data_in_1),
    .io_data_in_2(w8_a_io_data_in_2),
    .io_data_out(w8_a_io_data_out)
  );
  XOR32 w9_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w9_a_io_data_in_1),
    .io_data_in_2(w9_a_io_data_in_2),
    .io_data_out(w9_a_io_data_out)
  );
  XOR32 w10_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w10_a_io_data_in_1),
    .io_data_in_2(w10_a_io_data_in_2),
    .io_data_out(w10_a_io_data_out)
  );
  XOR32 w11_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w11_a_io_data_in_1),
    .io_data_in_2(w11_a_io_data_in_2),
    .io_data_out(w11_a_io_data_out)
  );
  ShiftRows data_c2_SR ( // @[ShiftRows.scala 14:20]
    .io_data_in(data_c2_SR_io_data_in),
    .io_data_out(data_c2_SR_io_data_out)
  );
  BS_MC data_c2_m ( // @[BS_MC.scala 72:19]
    .io_data_in(data_c2_m_io_data_in),
    .io_data_out(data_c2_m_io_data_out)
  );
  XOR128 round2_data_out_a ( // @[XOR32.scala 22:19]
    .io_data_in_1(round2_data_out_a_io_data_in_1),
    .io_data_in_2(round2_data_out_a_io_data_in_2),
    .io_data_out(round2_data_out_a_io_data_out)
  );
  G_func w12_g ( // @[G_func.scala 14:19]
    .io_data_in(w12_g_io_data_in),
    .io_rc_in(w12_g_io_rc_in),
    .io_data_out(w12_g_io_data_out)
  );
  XOR32 w12_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w12_a_io_data_in_1),
    .io_data_in_2(w12_a_io_data_in_2),
    .io_data_out(w12_a_io_data_out)
  );
  XOR32 w13_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w13_a_io_data_in_1),
    .io_data_in_2(w13_a_io_data_in_2),
    .io_data_out(w13_a_io_data_out)
  );
  XOR32 w14_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w14_a_io_data_in_1),
    .io_data_in_2(w14_a_io_data_in_2),
    .io_data_out(w14_a_io_data_out)
  );
  XOR32 w15_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w15_a_io_data_in_1),
    .io_data_in_2(w15_a_io_data_in_2),
    .io_data_out(w15_a_io_data_out)
  );
  ShiftRows data_c3_SR ( // @[ShiftRows.scala 14:20]
    .io_data_in(data_c3_SR_io_data_in),
    .io_data_out(data_c3_SR_io_data_out)
  );
  BS_MC data_c3_m ( // @[BS_MC.scala 72:19]
    .io_data_in(data_c3_m_io_data_in),
    .io_data_out(data_c3_m_io_data_out)
  );
  XOR128 round3_data_out_a ( // @[XOR32.scala 22:19]
    .io_data_in_1(round3_data_out_a_io_data_in_1),
    .io_data_in_2(round3_data_out_a_io_data_in_2),
    .io_data_out(round3_data_out_a_io_data_out)
  );
  G_func w16_g ( // @[G_func.scala 14:19]
    .io_data_in(w16_g_io_data_in),
    .io_rc_in(w16_g_io_rc_in),
    .io_data_out(w16_g_io_data_out)
  );
  XOR32 w16_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w16_a_io_data_in_1),
    .io_data_in_2(w16_a_io_data_in_2),
    .io_data_out(w16_a_io_data_out)
  );
  XOR32 w17_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w17_a_io_data_in_1),
    .io_data_in_2(w17_a_io_data_in_2),
    .io_data_out(w17_a_io_data_out)
  );
  XOR32 w18_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w18_a_io_data_in_1),
    .io_data_in_2(w18_a_io_data_in_2),
    .io_data_out(w18_a_io_data_out)
  );
  XOR32 w19_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w19_a_io_data_in_1),
    .io_data_in_2(w19_a_io_data_in_2),
    .io_data_out(w19_a_io_data_out)
  );
  ShiftRows data_c4_SR ( // @[ShiftRows.scala 14:20]
    .io_data_in(data_c4_SR_io_data_in),
    .io_data_out(data_c4_SR_io_data_out)
  );
  BS_MC data_c4_m ( // @[BS_MC.scala 72:19]
    .io_data_in(data_c4_m_io_data_in),
    .io_data_out(data_c4_m_io_data_out)
  );
  XOR128 round4_data_out_a ( // @[XOR32.scala 22:19]
    .io_data_in_1(round4_data_out_a_io_data_in_1),
    .io_data_in_2(round4_data_out_a_io_data_in_2),
    .io_data_out(round4_data_out_a_io_data_out)
  );
  G_func w20_g ( // @[G_func.scala 14:19]
    .io_data_in(w20_g_io_data_in),
    .io_rc_in(w20_g_io_rc_in),
    .io_data_out(w20_g_io_data_out)
  );
  XOR32 w20_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w20_a_io_data_in_1),
    .io_data_in_2(w20_a_io_data_in_2),
    .io_data_out(w20_a_io_data_out)
  );
  XOR32 w21_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w21_a_io_data_in_1),
    .io_data_in_2(w21_a_io_data_in_2),
    .io_data_out(w21_a_io_data_out)
  );
  XOR32 w22_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w22_a_io_data_in_1),
    .io_data_in_2(w22_a_io_data_in_2),
    .io_data_out(w22_a_io_data_out)
  );
  XOR32 w23_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w23_a_io_data_in_1),
    .io_data_in_2(w23_a_io_data_in_2),
    .io_data_out(w23_a_io_data_out)
  );
  ShiftRows data_c5_SR ( // @[ShiftRows.scala 14:20]
    .io_data_in(data_c5_SR_io_data_in),
    .io_data_out(data_c5_SR_io_data_out)
  );
  BS_MC data_c5_m ( // @[BS_MC.scala 72:19]
    .io_data_in(data_c5_m_io_data_in),
    .io_data_out(data_c5_m_io_data_out)
  );
  XOR128 round5_data_out_a ( // @[XOR32.scala 22:19]
    .io_data_in_1(round5_data_out_a_io_data_in_1),
    .io_data_in_2(round5_data_out_a_io_data_in_2),
    .io_data_out(round5_data_out_a_io_data_out)
  );
  G_func w24_g ( // @[G_func.scala 14:19]
    .io_data_in(w24_g_io_data_in),
    .io_rc_in(w24_g_io_rc_in),
    .io_data_out(w24_g_io_data_out)
  );
  XOR32 w24_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w24_a_io_data_in_1),
    .io_data_in_2(w24_a_io_data_in_2),
    .io_data_out(w24_a_io_data_out)
  );
  XOR32 w25_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w25_a_io_data_in_1),
    .io_data_in_2(w25_a_io_data_in_2),
    .io_data_out(w25_a_io_data_out)
  );
  XOR32 w26_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w26_a_io_data_in_1),
    .io_data_in_2(w26_a_io_data_in_2),
    .io_data_out(w26_a_io_data_out)
  );
  XOR32 w27_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w27_a_io_data_in_1),
    .io_data_in_2(w27_a_io_data_in_2),
    .io_data_out(w27_a_io_data_out)
  );
  ShiftRows data_c6_SR ( // @[ShiftRows.scala 14:20]
    .io_data_in(data_c6_SR_io_data_in),
    .io_data_out(data_c6_SR_io_data_out)
  );
  BS_MC data_c6_m ( // @[BS_MC.scala 72:19]
    .io_data_in(data_c6_m_io_data_in),
    .io_data_out(data_c6_m_io_data_out)
  );
  XOR128 round6_data_out_a ( // @[XOR32.scala 22:19]
    .io_data_in_1(round6_data_out_a_io_data_in_1),
    .io_data_in_2(round6_data_out_a_io_data_in_2),
    .io_data_out(round6_data_out_a_io_data_out)
  );
  G_func w28_g ( // @[G_func.scala 14:19]
    .io_data_in(w28_g_io_data_in),
    .io_rc_in(w28_g_io_rc_in),
    .io_data_out(w28_g_io_data_out)
  );
  XOR32 w28_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w28_a_io_data_in_1),
    .io_data_in_2(w28_a_io_data_in_2),
    .io_data_out(w28_a_io_data_out)
  );
  XOR32 w29_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w29_a_io_data_in_1),
    .io_data_in_2(w29_a_io_data_in_2),
    .io_data_out(w29_a_io_data_out)
  );
  XOR32 w30_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w30_a_io_data_in_1),
    .io_data_in_2(w30_a_io_data_in_2),
    .io_data_out(w30_a_io_data_out)
  );
  XOR32 w31_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w31_a_io_data_in_1),
    .io_data_in_2(w31_a_io_data_in_2),
    .io_data_out(w31_a_io_data_out)
  );
  ShiftRows data_c7_SR ( // @[ShiftRows.scala 14:20]
    .io_data_in(data_c7_SR_io_data_in),
    .io_data_out(data_c7_SR_io_data_out)
  );
  BS_MC data_c7_m ( // @[BS_MC.scala 72:19]
    .io_data_in(data_c7_m_io_data_in),
    .io_data_out(data_c7_m_io_data_out)
  );
  XOR128 round7_data_out_a ( // @[XOR32.scala 22:19]
    .io_data_in_1(round7_data_out_a_io_data_in_1),
    .io_data_in_2(round7_data_out_a_io_data_in_2),
    .io_data_out(round7_data_out_a_io_data_out)
  );
  G_func w32_g ( // @[G_func.scala 14:19]
    .io_data_in(w32_g_io_data_in),
    .io_rc_in(w32_g_io_rc_in),
    .io_data_out(w32_g_io_data_out)
  );
  XOR32 w32_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w32_a_io_data_in_1),
    .io_data_in_2(w32_a_io_data_in_2),
    .io_data_out(w32_a_io_data_out)
  );
  XOR32 w33_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w33_a_io_data_in_1),
    .io_data_in_2(w33_a_io_data_in_2),
    .io_data_out(w33_a_io_data_out)
  );
  XOR32 w34_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w34_a_io_data_in_1),
    .io_data_in_2(w34_a_io_data_in_2),
    .io_data_out(w34_a_io_data_out)
  );
  XOR32 w35_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w35_a_io_data_in_1),
    .io_data_in_2(w35_a_io_data_in_2),
    .io_data_out(w35_a_io_data_out)
  );
  ShiftRows data_c8_SR ( // @[ShiftRows.scala 14:20]
    .io_data_in(data_c8_SR_io_data_in),
    .io_data_out(data_c8_SR_io_data_out)
  );
  BS_MC data_c8_m ( // @[BS_MC.scala 72:19]
    .io_data_in(data_c8_m_io_data_in),
    .io_data_out(data_c8_m_io_data_out)
  );
  XOR128 round8_data_out_a ( // @[XOR32.scala 22:19]
    .io_data_in_1(round8_data_out_a_io_data_in_1),
    .io_data_in_2(round8_data_out_a_io_data_in_2),
    .io_data_out(round8_data_out_a_io_data_out)
  );
  G_func w36_g ( // @[G_func.scala 14:19]
    .io_data_in(w36_g_io_data_in),
    .io_rc_in(w36_g_io_rc_in),
    .io_data_out(w36_g_io_data_out)
  );
  XOR32 w36_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w36_a_io_data_in_1),
    .io_data_in_2(w36_a_io_data_in_2),
    .io_data_out(w36_a_io_data_out)
  );
  XOR32 w37_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w37_a_io_data_in_1),
    .io_data_in_2(w37_a_io_data_in_2),
    .io_data_out(w37_a_io_data_out)
  );
  XOR32 w38_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w38_a_io_data_in_1),
    .io_data_in_2(w38_a_io_data_in_2),
    .io_data_out(w38_a_io_data_out)
  );
  XOR32 w39_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w39_a_io_data_in_1),
    .io_data_in_2(w39_a_io_data_in_2),
    .io_data_out(w39_a_io_data_out)
  );
  ShiftRows data_c9_SR ( // @[ShiftRows.scala 14:20]
    .io_data_in(data_c9_SR_io_data_in),
    .io_data_out(data_c9_SR_io_data_out)
  );
  BS_MC data_c9_m ( // @[BS_MC.scala 72:19]
    .io_data_in(data_c9_m_io_data_in),
    .io_data_out(data_c9_m_io_data_out)
  );
  XOR128 round9_data_out_a ( // @[XOR32.scala 22:19]
    .io_data_in_1(round9_data_out_a_io_data_in_1),
    .io_data_in_2(round9_data_out_a_io_data_in_2),
    .io_data_out(round9_data_out_a_io_data_out)
  );
  G_func w40_g ( // @[G_func.scala 14:19]
    .io_data_in(w40_g_io_data_in),
    .io_rc_in(w40_g_io_rc_in),
    .io_data_out(w40_g_io_data_out)
  );
  XOR32 w40_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w40_a_io_data_in_1),
    .io_data_in_2(w40_a_io_data_in_2),
    .io_data_out(w40_a_io_data_out)
  );
  XOR32 w41_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w41_a_io_data_in_1),
    .io_data_in_2(w41_a_io_data_in_2),
    .io_data_out(w41_a_io_data_out)
  );
  XOR32 w42_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w42_a_io_data_in_1),
    .io_data_in_2(w42_a_io_data_in_2),
    .io_data_out(w42_a_io_data_out)
  );
  XOR32 w43_a ( // @[XOR32.scala 9:19]
    .io_data_in_1(w43_a_io_data_in_1),
    .io_data_in_2(w43_a_io_data_in_2),
    .io_data_out(w43_a_io_data_out)
  );
  ShiftRows data_c10_SR ( // @[ShiftRows.scala 14:20]
    .io_data_in(data_c10_SR_io_data_in),
    .io_data_out(data_c10_SR_io_data_out)
  );
  BS data_c10_m ( // @[BS_MC.scala 88:19]
    .io_data_in(data_c10_m_io_data_in),
    .io_data_out(data_c10_m_io_data_out)
  );
  XOR128 round10_data_out_a ( // @[XOR32.scala 22:19]
    .io_data_in_1(round10_data_out_a_io_data_in_1),
    .io_data_in_2(round10_data_out_a_io_data_in_2),
    .io_data_out(round10_data_out_a_io_data_out)
  );
  assign io_data_out = round10_data_out_a_io_data_out; // @[AES128.scala 226:30 AES128.scala 239:20]
  assign round0_data_out_a_io_data_in_1 = data_r0; // @[XOR32.scala 23:20]
  assign round0_data_out_a_io_data_in_2 = key_r0; // @[XOR32.scala 24:20]
  assign w4_g_io_data_in = key_r0[127:96]; // @[AES128.scala 29:28]
  assign w4_g_io_rc_in = 8'h1; // @[G_func.scala 16:16]
  assign w4_a_io_data_in_1 = w4_g_io_data_out; // @[XOR32.scala 10:20]
  assign w4_a_io_data_in_2 = key_r0[31:0]; // @[AES128.scala 29:60]
  assign w5_a_io_data_in_1 = w4_a_io_data_out; // @[AES128.scala 23:16 AES128.scala 29:6]
  assign w5_a_io_data_in_2 = key_r0[63:32]; // @[AES128.scala 30:25]
  assign w6_a_io_data_in_1 = w5_a_io_data_out; // @[AES128.scala 24:16 AES128.scala 30:6]
  assign w6_a_io_data_in_2 = key_r0[95:64]; // @[AES128.scala 31:25]
  assign w7_a_io_data_in_1 = w6_a_io_data_out; // @[AES128.scala 25:16 AES128.scala 31:6]
  assign w7_a_io_data_in_2 = key_r0[127:96]; // @[AES128.scala 32:25]
  assign data_c1_SR_io_data_in = round0_data_out_a_io_data_out; // @[AES128.scala 11:29 AES128.scala 19:19]
  assign data_c1_m_io_data_in = data_c1_SR_io_data_out; // @[BS_MC.scala 73:18]
  assign round1_data_out_a_io_data_in_1 = data_r1; // @[XOR32.scala 23:20]
  assign round1_data_out_a_io_data_in_2 = key_r1; // @[XOR32.scala 24:20]
  assign w8_g_io_data_in = key_r1[127:96]; // @[AES128.scala 51:28]
  assign w8_g_io_rc_in = 8'h2; // @[G_func.scala 16:16]
  assign w8_a_io_data_in_1 = w8_g_io_data_out; // @[XOR32.scala 10:20]
  assign w8_a_io_data_in_2 = key_r1[31:0]; // @[AES128.scala 51:60]
  assign w9_a_io_data_in_1 = w8_a_io_data_out; // @[AES128.scala 45:16 AES128.scala 51:6]
  assign w9_a_io_data_in_2 = key_r1[63:32]; // @[AES128.scala 52:25]
  assign w10_a_io_data_in_1 = w9_a_io_data_out; // @[AES128.scala 46:16 AES128.scala 52:6]
  assign w10_a_io_data_in_2 = key_r1[95:64]; // @[AES128.scala 53:26]
  assign w11_a_io_data_in_1 = w10_a_io_data_out; // @[AES128.scala 47:17 AES128.scala 53:7]
  assign w11_a_io_data_in_2 = key_r1[127:96]; // @[AES128.scala 54:27]
  assign data_c2_SR_io_data_in = round1_data_out_a_io_data_out; // @[AES128.scala 28:29 AES128.scala 41:19]
  assign data_c2_m_io_data_in = data_c2_SR_io_data_out; // @[BS_MC.scala 73:18]
  assign round2_data_out_a_io_data_in_1 = data_r2; // @[XOR32.scala 23:20]
  assign round2_data_out_a_io_data_in_2 = key_r2; // @[XOR32.scala 24:20]
  assign w12_g_io_data_in = key_r2[127:96]; // @[AES128.scala 73:29]
  assign w12_g_io_rc_in = 8'h4; // @[G_func.scala 16:16]
  assign w12_a_io_data_in_1 = w12_g_io_data_out; // @[XOR32.scala 10:20]
  assign w12_a_io_data_in_2 = key_r2[31:0]; // @[AES128.scala 73:61]
  assign w13_a_io_data_in_1 = w12_a_io_data_out; // @[AES128.scala 67:17 AES128.scala 73:7]
  assign w13_a_io_data_in_2 = key_r2[63:32]; // @[AES128.scala 74:27]
  assign w14_a_io_data_in_1 = w13_a_io_data_out; // @[AES128.scala 68:17 AES128.scala 74:7]
  assign w14_a_io_data_in_2 = key_r2[95:64]; // @[AES128.scala 75:27]
  assign w15_a_io_data_in_1 = w14_a_io_data_out; // @[AES128.scala 69:17 AES128.scala 75:7]
  assign w15_a_io_data_in_2 = key_r2[127:96]; // @[AES128.scala 76:27]
  assign data_c3_SR_io_data_in = round2_data_out_a_io_data_out; // @[AES128.scala 50:29 AES128.scala 63:19]
  assign data_c3_m_io_data_in = data_c3_SR_io_data_out; // @[BS_MC.scala 73:18]
  assign round3_data_out_a_io_data_in_1 = data_r3; // @[XOR32.scala 23:20]
  assign round3_data_out_a_io_data_in_2 = key_r3; // @[XOR32.scala 24:20]
  assign w16_g_io_data_in = key_r3[127:96]; // @[AES128.scala 95:29]
  assign w16_g_io_rc_in = 8'h8; // @[G_func.scala 16:16]
  assign w16_a_io_data_in_1 = w16_g_io_data_out; // @[XOR32.scala 10:20]
  assign w16_a_io_data_in_2 = key_r3[31:0]; // @[AES128.scala 95:61]
  assign w17_a_io_data_in_1 = w16_a_io_data_out; // @[AES128.scala 89:17 AES128.scala 95:7]
  assign w17_a_io_data_in_2 = key_r3[63:32]; // @[AES128.scala 96:27]
  assign w18_a_io_data_in_1 = w17_a_io_data_out; // @[AES128.scala 90:17 AES128.scala 96:7]
  assign w18_a_io_data_in_2 = key_r3[95:64]; // @[AES128.scala 97:27]
  assign w19_a_io_data_in_1 = w18_a_io_data_out; // @[AES128.scala 91:17 AES128.scala 97:7]
  assign w19_a_io_data_in_2 = key_r3[127:96]; // @[AES128.scala 98:27]
  assign data_c4_SR_io_data_in = round3_data_out_a_io_data_out; // @[AES128.scala 72:29 AES128.scala 85:19]
  assign data_c4_m_io_data_in = data_c4_SR_io_data_out; // @[BS_MC.scala 73:18]
  assign round4_data_out_a_io_data_in_1 = data_r4; // @[XOR32.scala 23:20]
  assign round4_data_out_a_io_data_in_2 = key_r4; // @[XOR32.scala 24:20]
  assign w20_g_io_data_in = key_r4[127:96]; // @[AES128.scala 117:29]
  assign w20_g_io_rc_in = 8'h10; // @[G_func.scala 16:16]
  assign w20_a_io_data_in_1 = w20_g_io_data_out; // @[XOR32.scala 10:20]
  assign w20_a_io_data_in_2 = key_r4[31:0]; // @[AES128.scala 117:61]
  assign w21_a_io_data_in_1 = w20_a_io_data_out; // @[AES128.scala 111:17 AES128.scala 117:7]
  assign w21_a_io_data_in_2 = key_r4[63:32]; // @[AES128.scala 118:27]
  assign w22_a_io_data_in_1 = w21_a_io_data_out; // @[AES128.scala 112:17 AES128.scala 118:7]
  assign w22_a_io_data_in_2 = key_r4[95:64]; // @[AES128.scala 119:27]
  assign w23_a_io_data_in_1 = w22_a_io_data_out; // @[AES128.scala 113:17 AES128.scala 119:7]
  assign w23_a_io_data_in_2 = key_r4[127:96]; // @[AES128.scala 120:27]
  assign data_c5_SR_io_data_in = round4_data_out_a_io_data_out; // @[AES128.scala 94:29 AES128.scala 107:19]
  assign data_c5_m_io_data_in = data_c5_SR_io_data_out; // @[BS_MC.scala 73:18]
  assign round5_data_out_a_io_data_in_1 = data_r5; // @[XOR32.scala 23:20]
  assign round5_data_out_a_io_data_in_2 = key_r5; // @[XOR32.scala 24:20]
  assign w24_g_io_data_in = key_r5[127:96]; // @[AES128.scala 139:29]
  assign w24_g_io_rc_in = 8'h20; // @[G_func.scala 16:16]
  assign w24_a_io_data_in_1 = w24_g_io_data_out; // @[XOR32.scala 10:20]
  assign w24_a_io_data_in_2 = key_r5[31:0]; // @[AES128.scala 139:61]
  assign w25_a_io_data_in_1 = w24_a_io_data_out; // @[AES128.scala 133:17 AES128.scala 139:7]
  assign w25_a_io_data_in_2 = key_r5[63:32]; // @[AES128.scala 140:27]
  assign w26_a_io_data_in_1 = w25_a_io_data_out; // @[AES128.scala 134:17 AES128.scala 140:7]
  assign w26_a_io_data_in_2 = key_r5[95:64]; // @[AES128.scala 141:27]
  assign w27_a_io_data_in_1 = w26_a_io_data_out; // @[AES128.scala 135:17 AES128.scala 141:7]
  assign w27_a_io_data_in_2 = key_r5[127:96]; // @[AES128.scala 142:27]
  assign data_c6_SR_io_data_in = round5_data_out_a_io_data_out; // @[AES128.scala 116:29 AES128.scala 129:19]
  assign data_c6_m_io_data_in = data_c6_SR_io_data_out; // @[BS_MC.scala 73:18]
  assign round6_data_out_a_io_data_in_1 = data_r6; // @[XOR32.scala 23:20]
  assign round6_data_out_a_io_data_in_2 = key_r6; // @[XOR32.scala 24:20]
  assign w28_g_io_data_in = key_r6[127:96]; // @[AES128.scala 161:29]
  assign w28_g_io_rc_in = 8'h40; // @[G_func.scala 16:16]
  assign w28_a_io_data_in_1 = w28_g_io_data_out; // @[XOR32.scala 10:20]
  assign w28_a_io_data_in_2 = key_r6[31:0]; // @[AES128.scala 161:61]
  assign w29_a_io_data_in_1 = w28_a_io_data_out; // @[AES128.scala 155:17 AES128.scala 161:7]
  assign w29_a_io_data_in_2 = key_r6[63:32]; // @[AES128.scala 162:27]
  assign w30_a_io_data_in_1 = w29_a_io_data_out; // @[AES128.scala 156:17 AES128.scala 162:7]
  assign w30_a_io_data_in_2 = key_r6[95:64]; // @[AES128.scala 163:27]
  assign w31_a_io_data_in_1 = w30_a_io_data_out; // @[AES128.scala 157:17 AES128.scala 163:7]
  assign w31_a_io_data_in_2 = key_r6[127:96]; // @[AES128.scala 164:27]
  assign data_c7_SR_io_data_in = round6_data_out_a_io_data_out; // @[AES128.scala 138:29 AES128.scala 151:19]
  assign data_c7_m_io_data_in = data_c7_SR_io_data_out; // @[BS_MC.scala 73:18]
  assign round7_data_out_a_io_data_in_1 = data_r7; // @[XOR32.scala 23:20]
  assign round7_data_out_a_io_data_in_2 = key_r7; // @[XOR32.scala 24:20]
  assign w32_g_io_data_in = key_r7[127:96]; // @[AES128.scala 183:29]
  assign w32_g_io_rc_in = 8'h80; // @[G_func.scala 16:16]
  assign w32_a_io_data_in_1 = w32_g_io_data_out; // @[XOR32.scala 10:20]
  assign w32_a_io_data_in_2 = key_r7[31:0]; // @[AES128.scala 183:61]
  assign w33_a_io_data_in_1 = w32_a_io_data_out; // @[AES128.scala 177:17 AES128.scala 183:7]
  assign w33_a_io_data_in_2 = key_r7[63:32]; // @[AES128.scala 184:27]
  assign w34_a_io_data_in_1 = w33_a_io_data_out; // @[AES128.scala 178:17 AES128.scala 184:7]
  assign w34_a_io_data_in_2 = key_r7[95:64]; // @[AES128.scala 185:27]
  assign w35_a_io_data_in_1 = w34_a_io_data_out; // @[AES128.scala 179:17 AES128.scala 185:7]
  assign w35_a_io_data_in_2 = key_r7[127:96]; // @[AES128.scala 186:27]
  assign data_c8_SR_io_data_in = round7_data_out_a_io_data_out; // @[AES128.scala 160:29 AES128.scala 173:19]
  assign data_c8_m_io_data_in = data_c8_SR_io_data_out; // @[BS_MC.scala 73:18]
  assign round8_data_out_a_io_data_in_1 = data_r8; // @[XOR32.scala 23:20]
  assign round8_data_out_a_io_data_in_2 = key_r8; // @[XOR32.scala 24:20]
  assign w36_g_io_data_in = key_r8[127:96]; // @[AES128.scala 205:29]
  assign w36_g_io_rc_in = 8'h1b; // @[G_func.scala 16:16]
  assign w36_a_io_data_in_1 = w36_g_io_data_out; // @[XOR32.scala 10:20]
  assign w36_a_io_data_in_2 = key_r8[31:0]; // @[AES128.scala 205:61]
  assign w37_a_io_data_in_1 = w36_a_io_data_out; // @[AES128.scala 199:17 AES128.scala 205:7]
  assign w37_a_io_data_in_2 = key_r8[63:32]; // @[AES128.scala 206:27]
  assign w38_a_io_data_in_1 = w37_a_io_data_out; // @[AES128.scala 200:17 AES128.scala 206:7]
  assign w38_a_io_data_in_2 = key_r8[95:64]; // @[AES128.scala 207:27]
  assign w39_a_io_data_in_1 = w38_a_io_data_out; // @[AES128.scala 201:17 AES128.scala 207:7]
  assign w39_a_io_data_in_2 = key_r8[127:96]; // @[AES128.scala 208:27]
  assign data_c9_SR_io_data_in = round8_data_out_a_io_data_out; // @[AES128.scala 182:29 AES128.scala 195:19]
  assign data_c9_m_io_data_in = data_c9_SR_io_data_out; // @[BS_MC.scala 73:18]
  assign round9_data_out_a_io_data_in_1 = data_r9; // @[XOR32.scala 23:20]
  assign round9_data_out_a_io_data_in_2 = key_r9; // @[XOR32.scala 24:20]
  assign w40_g_io_data_in = key_r9[127:96]; // @[AES128.scala 227:29]
  assign w40_g_io_rc_in = 8'h36; // @[G_func.scala 16:16]
  assign w40_a_io_data_in_1 = w40_g_io_data_out; // @[XOR32.scala 10:20]
  assign w40_a_io_data_in_2 = key_r9[31:0]; // @[AES128.scala 227:61]
  assign w41_a_io_data_in_1 = w40_a_io_data_out; // @[AES128.scala 221:17 AES128.scala 227:7]
  assign w41_a_io_data_in_2 = key_r9[63:32]; // @[AES128.scala 228:27]
  assign w42_a_io_data_in_1 = w41_a_io_data_out; // @[AES128.scala 222:17 AES128.scala 228:7]
  assign w42_a_io_data_in_2 = key_r9[95:64]; // @[AES128.scala 229:27]
  assign w43_a_io_data_in_1 = w42_a_io_data_out; // @[AES128.scala 223:17 AES128.scala 229:7]
  assign w43_a_io_data_in_2 = key_r9[127:96]; // @[AES128.scala 230:27]
  assign data_c10_SR_io_data_in = round9_data_out_a_io_data_out; // @[AES128.scala 204:29 AES128.scala 217:19]
  assign data_c10_m_io_data_in = data_c10_SR_io_data_out; // @[BS_MC.scala 89:18]
  assign round10_data_out_a_io_data_in_1 = data_r10; // @[XOR32.scala 23:20]
  assign round10_data_out_a_io_data_in_2 = key_r10; // @[XOR32.scala 24:20]
  always @(posedge clock) begin
    if (reset) begin // @[AES128.scala 12:23]
      data_r0 <= 128'h0; // @[AES128.scala 13:13]
    end else begin
      data_r0 <= io_data_in; // @[AES128.scala 16:13]
    end
    if (reset) begin // @[AES128.scala 12:23]
      key_r0 <= 128'h0; // @[AES128.scala 14:12]
    end else begin
      key_r0 <= io_key_in; // @[AES128.scala 17:12]
    end
    if (reset) begin // @[AES128.scala 34:23]
      data_r1 <= 128'h0; // @[AES128.scala 35:13]
    end else begin
      data_r1 <= data_c1; // @[AES128.scala 38:13]
    end
    if (reset) begin // @[AES128.scala 34:23]
      key_r1 <= 128'h0; // @[AES128.scala 36:12]
    end else begin
      key_r1 <= _key_r1_T; // @[AES128.scala 39:12]
    end
    if (reset) begin // @[AES128.scala 56:23]
      data_r2 <= 128'h0; // @[AES128.scala 57:13]
    end else begin
      data_r2 <= data_c2; // @[AES128.scala 60:13]
    end
    if (reset) begin // @[AES128.scala 56:23]
      key_r2 <= 128'h0; // @[AES128.scala 58:12]
    end else begin
      key_r2 <= _key_r2_T; // @[AES128.scala 61:12]
    end
    if (reset) begin // @[AES128.scala 78:23]
      data_r3 <= 128'h0; // @[AES128.scala 79:13]
    end else begin
      data_r3 <= data_c3; // @[AES128.scala 82:13]
    end
    if (reset) begin // @[AES128.scala 78:23]
      key_r3 <= 128'h0; // @[AES128.scala 80:12]
    end else begin
      key_r3 <= _key_r3_T; // @[AES128.scala 83:12]
    end
    if (reset) begin // @[AES128.scala 100:23]
      data_r4 <= 128'h0; // @[AES128.scala 101:13]
    end else begin
      data_r4 <= data_c4; // @[AES128.scala 104:13]
    end
    if (reset) begin // @[AES128.scala 100:23]
      key_r4 <= 128'h0; // @[AES128.scala 102:12]
    end else begin
      key_r4 <= _key_r4_T; // @[AES128.scala 105:12]
    end
    if (reset) begin // @[AES128.scala 122:23]
      data_r5 <= 128'h0; // @[AES128.scala 123:13]
    end else begin
      data_r5 <= data_c5; // @[AES128.scala 126:13]
    end
    if (reset) begin // @[AES128.scala 122:23]
      key_r5 <= 128'h0; // @[AES128.scala 124:12]
    end else begin
      key_r5 <= _key_r5_T; // @[AES128.scala 127:12]
    end
    if (reset) begin // @[AES128.scala 144:23]
      data_r6 <= 128'h0; // @[AES128.scala 145:13]
    end else begin
      data_r6 <= data_c6; // @[AES128.scala 148:13]
    end
    if (reset) begin // @[AES128.scala 144:23]
      key_r6 <= 128'h0; // @[AES128.scala 146:12]
    end else begin
      key_r6 <= _key_r6_T; // @[AES128.scala 149:12]
    end
    if (reset) begin // @[AES128.scala 166:23]
      data_r7 <= 128'h0; // @[AES128.scala 167:13]
    end else begin
      data_r7 <= data_c7; // @[AES128.scala 170:13]
    end
    if (reset) begin // @[AES128.scala 166:23]
      key_r7 <= 128'h0; // @[AES128.scala 168:12]
    end else begin
      key_r7 <= _key_r7_T; // @[AES128.scala 171:12]
    end
    if (reset) begin // @[AES128.scala 188:23]
      data_r8 <= 128'h0; // @[AES128.scala 189:13]
    end else begin
      data_r8 <= data_c8; // @[AES128.scala 192:13]
    end
    if (reset) begin // @[AES128.scala 188:23]
      key_r8 <= 128'h0; // @[AES128.scala 190:12]
    end else begin
      key_r8 <= _key_r8_T; // @[AES128.scala 193:12]
    end
    if (reset) begin // @[AES128.scala 210:23]
      data_r9 <= 128'h0; // @[AES128.scala 211:13]
    end else begin
      data_r9 <= data_c9; // @[AES128.scala 214:13]
    end
    if (reset) begin // @[AES128.scala 210:23]
      key_r9 <= 128'h0; // @[AES128.scala 212:12]
    end else begin
      key_r9 <= _key_r9_T; // @[AES128.scala 215:12]
    end
    if (reset) begin // @[AES128.scala 232:23]
      data_r10 <= 128'h0; // @[AES128.scala 233:14]
    end else begin
      data_r10 <= data_c10; // @[AES128.scala 236:14]
    end
    if (reset) begin // @[AES128.scala 232:23]
      key_r10 <= 128'h0; // @[AES128.scala 234:13]
    end else begin
      key_r10 <= _key_r10_T; // @[AES128.scala 237:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  data_r0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  key_r0 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  data_r1 = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  key_r1 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  data_r2 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  key_r2 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  data_r3 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  key_r3 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  data_r4 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  key_r4 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  data_r5 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  key_r5 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  data_r6 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  key_r6 = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  data_r7 = _RAND_14[127:0];
  _RAND_15 = {4{`RANDOM}};
  key_r7 = _RAND_15[127:0];
  _RAND_16 = {4{`RANDOM}};
  data_r8 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  key_r8 = _RAND_17[127:0];
  _RAND_18 = {4{`RANDOM}};
  data_r9 = _RAND_18[127:0];
  _RAND_19 = {4{`RANDOM}};
  key_r9 = _RAND_19[127:0];
  _RAND_20 = {4{`RANDOM}};
  data_r10 = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  key_r10 = _RAND_21[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
